C2837611|T037|S32.048B|ICD10CM|OTHER FRACTURE OF FOURTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF FOURTH LUMBAR VERTEBRA, INIT FOR OPN FX
C2837610|T037|S32.048A|ICD10CM|OTHER FRACTURE OF FOURTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF FOURTH LUMBAR VERTEBRA, INIT FOR CLOS FX
C2888721|T047|L97.509|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF UNSPECIFIED FOOT WITH UNSPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OTH PRT UNSP FOOT W UNSP SEVERITY
C4509313|T047|L97.508|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF UNSPECIFIED FOOT WITH OTHER SPECIFIED SEVERITY|NON-PRS CHRONIC ULCER OTH PRT UNSP FOOT WITH OTH SEVERITY
C4268080|T047|E11.3391|ICD10CM|TYPE 2 DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|TYPE 2 DIAB WITH MOD NONP RTNOP WITHOUT MACULAR EDEMA, R EYE
C4268082|T047|E11.3393|ICD10CM|TYPE 2 DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|TYPE 2 DIAB WITH MOD NONP RTNOP WITHOUT MACULAR EDEMA, BI
C4268081|T047|E11.3392|ICD10CM|TYPE 2 DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|TYPE 2 DIAB WITH MOD NONP RTNOP WITHOUT MACULAR EDEMA, L EYE
C2888719|T047|L97.503|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF UNSPECIFIED FOOT WITH NECROSIS OF MUSCLE|NON-PRS CHRONIC ULCER OTH PRT UNSP FOOT W NECROSIS OF MUSCLE
C2888718|T047|L97.502|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF UNSPECIFIED FOOT WITH FAT LAYER EXPOSED|NON-PRS CHRONIC ULCER OTH PRT UNSP FOOT W FAT LAYER EXPOSED
C2888717|T047|L97.501|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF UNSPECIFIED FOOT LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHR ULCER OTH PRT UNSP FOOT LIMITED TO BRKDWN SKIN
C4268083|T047|E11.3399|ICD10CM|TYPE 2 DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|TYPE 2 DIAB WITH MOD NONP RTNOP WITHOUT MACULAR EDEMA, UNSP
C4509312|T047|L97.506|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF UNSPECIFIED FOOT WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OTH PRT UNSP FT W BNE INVL W/O EVD OF NECR
C4509311|T047|L97.505|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF UNSPECIFIED FOOT WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OTH PRT UNSP FT W MSL INVL W/O EVD OF NECR
C2888720|T047|L97.504|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF UNSPECIFIED FOOT WITH NECROSIS OF BONE|NON-PRS CHRONIC ULCER OTH PRT UNSP FOOT W NECROSIS OF BONE
C2976979|T046|I82.409|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF UNSPECIFIED LOWER EXTREMITY|ACUTE EMBOLISM AND THOMBOS UNSP DEEP VN UNSP LOWER EXTREMITY
C2976978|T046|I82.403|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF LOWER EXTREMITY, BILATERAL|ACUTE EMBOLISM AND THOMBOS UNSP DEEP VEINS OF LOW EXTRM, BI
C2976977|T046|I82.402|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF LEFT LOWER EXTREMITY|ACUTE EMBOLISM AND THOMBOS UNSP DEEP VEINS OF L LOW EXTREM
C2976976|T046|I82.401|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF RIGHT LOWER EXTREMITY|ACUTE EMBOLISM AND THOMBOS UNSP DEEP VEINS OF R LOW EXTREM
C2855885|T037|S68.115S|ICD10CM|COMPLETE TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF LEFT RING FINGER, SEQUELA|COMPLETE TRAUMATIC MCP AMPUTATION OF L RNG FNGR, SEQUELA
C0220992|T047|E70.41|ICD10CM|HISTIDINEMIA|HISTIDINEMIA
C0268512|T047|E70.40|ICD10CM|DISORDERS OF HISTIDINE METABOLISM, UNSPECIFIED|DISORDERS OF HISTIDINE METABOLISM, UNSPECIFIED
C0238286|T047|E75.11|ICD10CM|MUCOLIPIDOSIS IV|MUCOLIPIDOSIS IV
C0017083|T047|E75.10|ICD10CM|UNSPECIFIED GANGLIOSIDOSIS|UNSPECIFIED GANGLIOSIDOSIS
C2874234|T047|E70.49|ICD10CM|OTHER DISORDERS OF HISTIDINE METABOLISM|OTHER DISORDERS OF HISTIDINE METABOLISM
C0795951|T047||ICD10CM|OTHER GANGLIOSIDOSIS
C2833927|T037|S14.123A|ICD10CM|CENTRAL CORD SYNDROME AT C3 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|CENTRAL CORD SYNDROME AT C3, INIT
C2874194|T047|E26.09|ICD10CM|OTHER PRIMARY HYPERALDOSTERONISM|OTHER PRIMARY HYPERALDOSTERONISM
C2831496|T037|S02.412S|ICD10CM|LEFORT II FRACTURE, SEQUELA|LEFORT II FRACTURE, SEQUELA
C2831491|T037|S02.412A|ICD10CM|LEFORT II FRACTURE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|LEFORT II FRACTURE, INITIAL ENCOUNTER FOR CLOSED FRACTURE
C2831492|T037|S02.412B|ICD10CM|LEFORT II FRACTURE, INITIAL ENCOUNTER FOR OPEN FRACTURE|LEFORT II FRACTURE, INITIAL ENCOUNTER FOR OPEN FRACTURE
C2882664|T047|I69.941|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING RIGHT DOMINANT SIDE|MONOPLG LOW LMB FOL UNSP CEREBVASC DIS AFF RIGHT DOM SIDE
C2878923|T037|T44.7X2S|ICD10CM|POISONING BY BETA-ADRENORECEPTOR ANTAGONISTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY BETA-ADRENOCPT ANTAGONISTS, SELF-HARM, SEQUELA
C2858628|T037|S72.436B|ICD10CM|NONDISPLACED FRACTURE OF MEDIAL CONDYLE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF MED CONDYLE OF UNSP FEMR, 7THB
C0838550|T047|M46.88|ICD10CM|OTHER SPECIFIED INFLAMMATORY SPONDYLOPATHIES, SACRAL AND SACROCOCCYGEAL REGION|OTH INFLAMMATORY SPONDYLOPATHIES, SACR/SACROCYGL REGION
C2883610|T037|T50.3X2A|ICD10CM|POISONING BY ELECTROLYTIC, CALORIC AND WATER-BALANCE AGENTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY ELECTROLYTIC/CALORIC/WTR-BAL AGNT, SELF-HARM, INIT
C2883057|T047|I80.13|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF FEMORAL VEIN, BILATERAL|PHLEBITIS AND THROMBOPHLEBITIS OF FEMORAL VEIN, BILATERAL
C0838551|T047|M46.89|ICD10AM|OTHER SPECIFIED INFLAMMATORY SPONDYLOPATHIES, MULTIPLE SITES IN SPINE|OTHER SPECIFIED INFLAMMATORY SPONDYLOPATHIES, SITE UNSPECIFIED
C2873872|T047|E05.31|ICD10CM|THYROTOXICOSIS FROM ECTOPIC THYROID TISSUE WITH THYROTOXIC CRISIS OR STORM|THYROTXCOSIS FROM ECTOPIC THYROID TISSUE W THYROTOXIC CRISIS
C2883056|T047|I80.12|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF LEFT FEMORAL VEIN|PHLEBITIS AND THROMBOPHLEBITIS OF LEFT FEMORAL VEIN
C4269585|T037|S02.82XS|ICD10CM|FRACTURE OF OTHER SPECIFIED SKULL AND FACIAL BONES, LEFT SIDE, SEQUELA|FRACTURE OF OTH SKULL AND FACIAL BONES, LEFT SIDE, SEQUELA
C2883612|T037|T50.3X2S|ICD10CM|POISONING BY ELECTROLYTIC, CALORIC AND WATER-BALANCE AGENTS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY ELECTROLYTIC/CALORIC/WTR-BAL AGNT, SLF-HRM, SEQUELA
C2883055|T047|I80.11|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF RIGHT FEMORAL VEIN|PHLEBITIS AND THROMBOPHLEBITIS OF RIGHT FEMORAL VEIN
C2882667|T047|I69.944|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING LEFT NON-DOMINANT SIDE|MONOPLG LOW LMB FOL UNSP CEREBVASC DIS AFF LEFT NONDOM SIDE
C2883054|T047|I80.10|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF UNSPECIFIED FEMORAL VEIN|PHLEBITIS AND THROMBOPHLEBITIS OF UNSPECIFIED FEMORAL VEIN
C4267963|T047|E09.3312|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|DRUG/CHEM DIAB WITH MOD NONP RTNOP WITH MACULAR EDEMA, L EYE
C4267964|T047|E09.3313|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|DRUG/CHEM DIAB WITH MOD NONP RTNOP WITH MACULAR EDEMA, BI
C4267962|T047|E09.3311|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|DRUG/CHEM DIAB WITH MOD NONP RTNOP WITH MACULAR EDEMA, R EYE
C2837720|T037|S32.129A|ICD10CM|UNSPECIFIED ZONE II FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP ZONE II FRACTURE OF SACRUM, INIT FOR CLOS FX
C2860007|T037|S78.119S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN UNSPECIFIED HIP AND KNEE, SEQUELA|COMPLETE TRAUM AMP AT LEVEL BETW UNSP HIP AND KNEE, SEQUELA
C4267965|T047|E09.3319|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|DRUG/CHEM DIAB WITH MOD NONP RTNOP WITH MACULAR EDEMA, UNSP
C0838544|T047|M46.82|ICD10CM|OTHER SPECIFIED INFLAMMATORY SPONDYLOPATHIES, CERVICAL REGION|OTH INFLAMMATORY SPONDYLOPATHIES, CERVICAL REGION
C2901004|T046|M84.453A|ICD10CM|PATHOLOGICAL FRACTURE, UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, UNSP FEMUR, INIT ENCNTR FOR FRACTURE
C2860005|T037|S78.119A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN UNSPECIFIED HIP AND KNEE, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMP AT LEVEL BETW UNSP HIP AND KNEE, INIT
C2860006|T037|S78.119D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN UNSPECIFIED HIP AND KNEE, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMP AT LEVEL BETW UNSP HIP AND KNEE, SUBS
C2902064|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, RIGHT TIBIA
C2902065|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, LEFT TIBIA
C2902066|T046|M87.263|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED TIBIA|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED TIBIA
C2902067|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, RIGHT FIBULA
C2902068|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, LEFT FIBULA
C2902069|T046|M87.266|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED FIBULA|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED FIBULA
C2877097|T037|T38.4X2A|ICD10CM|POISONING BY ORAL CONTRACEPTIVES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ORAL CONTRACEPTIVES, SELF-HARM, INIT
C0838549|T047|M46.87|ICD10CM|OTHER SPECIFIED INFLAMMATORY SPONDYLOPATHIES, LUMBOSACRAL REGION|OTH INFLAMMATORY SPONDYLOPATHIES, LUMBOSACRAL REGION
C2882078|T047|I12.0|ICD10CM|HYPERTENSIVE CHRONIC KIDNEY DISEASE WITH STAGE 5 CHRONIC KIDNEY DISEASE OR END STAGE RENAL DISEASE|HYP CHR KIDNEY DISEASE W STAGE 5 CHR KIDNEY DISEASE OR ESRD
C3695318|T047||ICD10CM|HYPERTENSIVE CHRONIC KIDNEY DISEASE WITH STAGE 1 THROUGH STAGE 4 CHRONIC KIDNEY DISEASE, OR UNSPECIFIED CHRONIC KIDNEY DISEASE
C2845912|T191|C69.41|ICD10CM|MALIGNANT NEOPLASM OF RIGHT CILIARY BODY|MALIGNANT NEOPLASM OF RIGHT CILIARY BODY
C2845911|T191|C69.40|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED CILIARY BODY|MALIGNANT NEOPLASM OF UNSPECIFIED CILIARY BODY
C2845913|T191|C69.42|ICD10CM|MALIGNANT NEOPLASM OF LEFT CILIARY BODY|MALIGNANT NEOPLASM OF LEFT CILIARY BODY
C2833628|T037|S12.651A|ICD10CM|OTHER TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH TRAUM NONDISP SPONDYLOLYSIS OF 7TH CERVCAL VERT, INIT
C2889420|T047|M06.229|ICD10CM|RHEUMATOID BURSITIS, UNSPECIFIED ELBOW|RHEUMATOID BURSITIS, UNSPECIFIED ELBOW
C2833629|T037|S12.651B|ICD10CM|OTHER TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH TRAUM NONDISP SPONDYLOLYSIS OF 7TH CERVCAL VERT, 7THB
C2858527|T037|S72.426C|ICD10CM|NONDISPLACED FRACTURE OF LATERAL CONDYLE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF LATERAL CONDYLE OF UNSP FEMR, 7THC
C2858526|T037|S72.426B|ICD10CM|NONDISPLACED FRACTURE OF LATERAL CONDYLE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF LATERAL CONDYLE OF UNSP FEMR, 7THB
C2858525|T037|S72.426A|ICD10CM|NONDISPLACED FRACTURE OF LATERAL CONDYLE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF LATERAL CONDYLE OF UNSP FEMUR, INIT
C2880026|T037|T48.3X2S|ICD10CM|POISONING BY ANTITUSSIVES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ANTITUSSIVES, INTENTIONAL SELF-HARM, SEQUELA
C2889419|T047|M06.222|ICD10CM|RHEUMATOID BURSITIS, LEFT ELBOW|RHEUMATOID BURSITIS, LEFT ELBOW
C2889418|T047|M06.221|ICD10CM|RHEUMATOID BURSITIS, RIGHT ELBOW|RHEUMATOID BURSITIS, RIGHT ELBOW
C2888026|T046|K94.09|ICD10CM|OTHER COMPLICATIONS OF COLOSTOMY|OTHER COMPLICATIONS OF COLOSTOMY
C0078918|T019|E70.329|ICD10CM|OCULOCUTANEOUS ALBINISM, UNSPECIFIED|OCULOCUTANEOUS ALBINISM, UNSPECIFIED
C2936910|T047|E70.328|ICD10CM|OTHER OCULOCUTANEOUS ALBINISM|CROSS SYNDROME
C2888025|T046|K94.01|ICD10CM|COLOSTOMY HEMORRHAGE|COLOSTOMY HEMORRHAGE
C2888024|T046|K94.00|ICD10CM|COLOSTOMY COMPLICATION, UNSPECIFIED|COLOSTOMY COMPLICATION, UNSPECIFIED
C2106483|T046|K94.03|ICD10CM|COLOSTOMY MALFUNCTION|MECHANICAL COMPLICATION OF COLOSTOMY
C0854424|T046|K94.02|ICD10CM|COLOSTOMY INFECTION|COLOSTOMY INFECTION
C2890080|T037|T82.534A|ICD10CM|LEAKAGE OF INFUSION CATHETER, INITIAL ENCOUNTER|LEAKAGE OF INFUSION CATHETER, INITIAL ENCOUNTER
C0268495|T047|E70.321|ICD10CM|TYROSINASE POSITIVE OCULOCUTANEOUS ALBINISM|OCULOCUTANEOUS ALBINISM TY-POS
C0268494|T047|E70.320|ICD10CM|TYROSINASE NEGATIVE OCULOCUTANEOUS ALBINISM|OCULOCUTANEOUS ALBINISM TY-NEG
C2832368|T037|S06.375S|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF CEREBELLUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, SEQUELA|CONTUS/LAC/HEM CRBLM W LOC >24 HR W RET CONSC LEV, SEQUELA
C2882101|T047|I21.11|ICD10CM|ST ELEVATION (STEMI) MYOCARDIAL INFARCTION INVOLVING RIGHT CORONARY ARTERY|STEMI INVOLVING RIGHT CORONARY ARTERY
C2889445|T046|M06.322|ICD10CM|RHEUMATOID NODULE, LEFT ELBOW|RHEUMATOID NODULE, LEFT ELBOW
C2889444|T046|M06.321|ICD10CM|RHEUMATOID NODULE, RIGHT ELBOW|RHEUMATOID NODULE, RIGHT ELBOW
C2832366|T037|S06.375A|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF CEREBELLUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, INITIAL ENCOUNTER|CONTUS/LAC/HEM CRBLM W LOC >24 HR W RET CONSC LEV, INIT
C2889446|T046|M06.329|ICD10CM|RHEUMATOID NODULE, UNSPECIFIED ELBOW|RHEUMATOID NODULE, UNSPECIFIED ELBOW
C2883206|T037|T48.6X2S|ICD10CM|POISONING BY ANTIASTHMATICS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ANTIASTHMATICS, INTENTIONAL SELF-HARM, SEQUELA
C2879848|T037|T47.7X2S|ICD10CM|POISONING BY EMETICS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY EMETICS, INTENTIONAL SELF-HARM, SEQUELA
C2902855|T047|N00.9|ICD10CM|ACUTE NEPHRITIC SYNDROME WITH UNSPECIFIED MORPHOLOGIC CHANGES|ACUTE NEPHRITIC SYNDROME WITH UNSP MORPHOLOGIC CHANGES
C2883204|T037|T48.6X2A|ICD10CM|POISONING BY ANTIASTHMATICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ANTIASTHMATICS, INTENTIONAL SELF-HARM, INIT
C3665551|T191||ICD10CM|MALIGNANT NEOPLASM OF NASOPHARYNX, UNSPECIFIED
C0349038|T191|C11.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF NASOPHARYNX|BOESARTIGE NEUBILDUNG: NASOPHARYNX, MEHRERE TEILBEREICHE UEBERLAPPEND
C2833850|T191|C11.3|ICD10CM|MALIGNANT NEOPLASM OF ANTERIOR WALL OF NASOPHARYNX|MALIGNANT NEOPLASM OF POSTERIOR MARGIN OF NASAL SEPTUM
C0345658|T191|C11.2|ICD10CM|MALIGNANT NEOPLASM OF LATERAL WALL OF NASOPHARYNX|MALIGNANT NEOPLASM OF OPENING OF AUDITORY TUBE
C0345653|T191|C11.1|ICD10CM|MALIGNANT NEOPLASM OF POSTERIOR WALL OF NASOPHARYNX|MALIGNANT NEOPLASM OF ADENOID
C0153393|T191|C11.0|DMDICD10|MALIGNANT NEOPLASM OF SUPERIOR WALL OF NASOPHARYNX|BOESARTIGE NEUBILDUNG: OBERE WAND DES NASOPHARYNX
C2887754|T047|K50.011|ICD10CM|CROHN'S DISEASE OF SMALL INTESTINE WITH RECTAL BLEEDING|CROHN'S DISEASE OF SMALL INTESTINE WITH RECTAL BLEEDING
C2887756|T047|K50.013|ICD10CM|CROHN'S DISEASE OF SMALL INTESTINE WITH FISTULA|CROHN'S DISEASE OF SMALL INTESTINE WITH FISTULA
C2887755|T047|K50.012|ICD10CM|CROHN'S DISEASE OF SMALL INTESTINE WITH INTESTINAL OBSTRUCTION|CROHN'S DISEASE OF SMALL INTESTINE W INTESTINAL OBSTRUCTION
C2887757|T047|K50.014|ICD10CM|CROHN'S DISEASE OF SMALL INTESTINE WITH ABSCESS|CROHN'S DISEASE OF SMALL INTESTINE WITH ABSCESS
C2861666|T191|D03.11|ICD10CM|MELANOMA IN SITU OF RIGHT EYELID, INCLUDING CANTHUS|MELANOMA IN SITU OF RIGHT EYELID, INCLUDING CANTHUS
C2861665|T191|D03.10|ICD10CM|MELANOMA IN SITU OF UNSPECIFIED EYELID, INCLUDING CANTHUS|MELANOMA IN SITU OF UNSPECIFIED EYELID, INCLUDING CANTHUS
C2861667|T191|D03.12|ICD10CM|MELANOMA IN SITU OF LEFT EYELID, INCLUDING CANTHUS|MELANOMA IN SITU OF LEFT EYELID, INCLUDING CANTHUS
C2837691|T037|S32.119B|ICD10CM|UNSPECIFIED ZONE I FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP ZONE I FRACTURE OF SACRUM, INIT FOR OPN FX
C2837690|T037|S32.119A|ICD10CM|UNSPECIFIED ZONE I FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP ZONE I FRACTURE OF SACRUM, INIT FOR CLOS FX
C0154195|T047|E21.4|DMDICD10|OTHER SPECIFIED DISORDERS OF PARATHYROID GLAND|SONSTIGE NAEHER BEZEICHNETE KRANKHEITEN DER NEBENSCHILDDRUESE
C0030517|T047|E21.5|DMDICD10|DISORDER OF PARATHYROID GLAND, UNSPECIFIED|KRANKHEIT DER NEBENSCHILDDRUESE, NICHT NAEHER BEZEICHNET
C0348455|T047|E21.2|DMDICD10|OTHER HYPERPARATHYROIDISM|SONSTIGER HYPERPARATHYREOIDISMUS
C0020502|T047|E21.3|DMDICD10|HYPERPARATHYROIDISM, UNSPECIFIED|HYPERPARATHYREOIDISMUS, NICHT NAEHER BEZEICHNET
C2874186|T047|E21.0|ICD10CM|PRIMARY HYPERPARATHYROIDISM|OSTEITIS FIBROSA CYSTICA GENERALISATA [VON RECKLINGHAUSEN'S DISEASE OF BONE]
C0494305|T047|E21.1|DMDICD10|SECONDARY HYPERPARATHYROIDISM, NOT ELSEWHERE CLASSIFIED|SEKUNDAERER HYPERPARATHYREOIDISMUS, ANDERENORTS NICHT KLASSIFIZIERT
C0348487|T047|E74.8|DMDICD10|OTHER SPECIFIED DISORDERS OF CARBOHYDRATE METABOLISM|SONSTIGE NAEHER BEZEICHNETE STOERUNGEN DES KOHLENHYDRATSTOFFWECHSELS
C0149670|T047|E74.9|DMDICD10|DISORDER OF CARBOHYDRATE METABOLISM, UNSPECIFIED|STOERUNG DES KOHLENHYDRATSTOFFWECHSELS, NICHT NAEHER BEZEICHNET
C4269389|T037|S02.40BS|ICD10CM|MALAR FRACTURE, LEFT SIDE, SEQUELA|MALAR FRACTURE, LEFT SIDE, SEQUELA
C2888417|T047|L89.302|ICD10CM|PRESSURE ULCER OF UNSPECIFIED BUTTOCK, STAGE 2|PRESSURE ULCER OF UNSPECIFIED BUTTOCK, STAGE 2
C2888420|T047|L89.303|ICD10CM|PRESSURE ULCER OF UNSPECIFIED BUTTOCK, STAGE 3|PRESSURE ULCER OF UNSPECIFIED BUTTOCK, STAGE 3
C2888411|T047|L89.300|ICD10CM|PRESSURE ULCER OF UNSPECIFIED BUTTOCK, UNSTAGEABLE|PRESSURE ULCER OF UNSPECIFIED BUTTOCK, UNSTAGEABLE
C2888414|T047|L89.301|ICD10CM|PRESSURE ULCER OF UNSPECIFIED BUTTOCK, STAGE 1|PRESSURE ULCER OF UNSPECIFIED BUTTOCK, STAGE 1
C2888423|T047|L89.304|ICD10CM|PRESSURE ULCER OF UNSPECIFIED BUTTOCK, STAGE 4|PRESSURE ULCER OF UNSPECIFIED BUTTOCK, STAGE 4
C4269384|T037|S02.40BA|ICD10CM|MALAR FRACTURE, LEFT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|MALAR FRACTURE, LEFT SIDE, INIT
C4269385|T037|S02.40BB|ICD10CM|MALAR FRACTURE, LEFT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|MALAR FRACTURE, LEFT SIDE, 7THB
C2888426|T047|L89.309|ICD10CM|PRESSURE ULCER OF UNSPECIFIED BUTTOCK, UNSPECIFIED STAGE|PRESSURE ULCER OF UNSPECIFIED BUTTOCK, UNSPECIFIED STAGE
C2838035|T037|S32.415A|ICD10CM|NONDISPLACED FRACTURE OF ANTERIOR WALL OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF ANTERIOR WALL OF LEFT ACETABULUM, INIT
C2838230|T037|S32.462B|ICD10CM|DISPLACED ASSOCIATED TRANSVERSE-POSTERIOR FRACTURE OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISPLACED ASSOC TRANSV/POST FX LEFT ACETAB, INIT FOR OPN FX
C2838229|T037|S32.462A|ICD10CM|DISPLACED ASSOCIATED TRANSVERSE-POSTERIOR FRACTURE OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED ASSOCIATED TRANSV/POST FX LEFT ACETABULUM, INIT
C2838036|T037|S32.415B|ICD10CM|NONDISPLACED FRACTURE OF ANTERIOR WALL OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP FX OF ANTERIOR WALL OF LEFT ACETAB, INIT FOR OPN FX
C2882773|T047|I70.338|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF OTHER PART OF LOWER LEG|ATHSCL UNSP TYPE BYPASS OF RIGHT LEG W ULCER OTH PRT LOW LEG
C2837729|T037|S32.130A|ICD10CM|NONDISPLACED ZONE III FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED ZONE III FRACTURE OF SACRUM, INIT FOR CLOS FX
C2882774|T047|I70.339|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF UNSPECIFIED SITE|ATHSCL UNSP TYPE BYPASS OF RIGHT LEG W ULCER OF UNSP SITE
C2869764|T037|S98.019D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED FOOT AT ANKLE LEVEL, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMP OF UNSP FOOT AT ANKLE LEVEL, SUBS
C2837983|T191|C40.91|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED BONES AND ARTICULAR CARTILAGE OF RIGHT LIMB|MALIG NEOPLASM OF UNSP BONES AND ARTIC CARTLG OF RIGHT LIMB
C2837982|T191|C40.90|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED BONES AND ARTICULAR CARTILAGE OF UNSPECIFIED LIMB|MALIG NEOPLASM OF UNSP BONES AND ARTIC CARTLG OF UNSP LIMB
C2837984|T191|C40.92|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED BONES AND ARTICULAR CARTILAGE OF LEFT LIMB|MALIG NEOPLASM OF UNSP BONES AND ARTIC CARTLG OF LEFT LIMB
C2900441|T047||ICD10CM|ARTHRITIS DUE TO LYME DISEASE
C2860193|T037|S79.132A|ICD10CM|SALTER-HARRIS TYPE III PHYSEAL FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SLTR-HARIS TYPE III PHYSEAL FX LOWER END OF LEFT FEMUR, INIT
C2893648|T047|M12.061|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], RIGHT KNEE|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], RIGHT KNEE
C2889467|T047|M06.811|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, RIGHT SHOULDER|OTHER SPECIFIED RHEUMATOID ARTHRITIS, RIGHT SHOULDER
C2889468|T047|M06.812|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, LEFT SHOULDER|OTHER SPECIFIED RHEUMATOID ARTHRITIS, LEFT SHOULDER
C2902443|T047|M90.559|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, UNSPECIFIED THIGH|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, UNSP THIGH
C4270344|T046|T83.593A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO OTHER URINARY STENTS, INITIAL ENCOUNTER|I/I REACT D/T OTHER URINARY STENTS, INITIAL ENCOUNTER
C2848402|T037|S58.021A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT ELBOW LEVEL, RIGHT ARM, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION AT ELBOW LEVEL, RIGHT ARM, INIT
C2902442|T047|M90.552|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, LEFT THIGH|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, LEFT THIGH
C2889469|T047|M06.819|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, UNSPECIFIED SHOULDER|OTHER SPECIFIED RHEUMATOID ARTHRITIS, UNSPECIFIED SHOULDER
C2911632|T047|B37.7|ICD10CM|CANDIDAL SEPSIS|CANDIDAL SEPSIS
C2911629|T047|B37.1|ICD10CM|PULMONARY CANDIDIASIS|CANDIDAL BRONCHITIS
C2848404|T037|S58.021S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT ELBOW LEVEL, RIGHT ARM, SEQUELA|PARTIAL TRAUMATIC AMP AT ELBOW LEVEL, RIGHT ARM, SEQUELA
C2889939|T037|T82.331A|ICD10CM|LEAKAGE OF CAROTID ARTERIAL GRAFT (BYPASS), INITIAL ENCOUNTER|LEAKAGE OF CAROTID ARTERIAL GRAFT (BYPASS), INIT ENCNTR
C2874292|T047|E78.70|ICD10CM|DISORDER OF BILE ACID AND CHOLESTEROL METABOLISM, UNSPECIFIED|DISORDER OF BILE ACID AND CHOLESTEROL METABOLISM, UNSP
C2832317|T037|S06.363A|ICD10CM|TRAUMATIC HEMORRHAGE OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF 1 HOURS TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|TRAUM HEMOR CEREB, W LOC OF 1-5 HRS 59 MINUTES, INIT
C2874293|T047|E78.79|ICD10CM|OTHER DISORDERS OF BILE ACID AND CHOLESTEROL METABOLISM|OTHER DISORDERS OF BILE ACID AND CHOLESTEROL METABOLISM
C2893650|T047|M12.069|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], UNSPECIFIED KNEE|CHRONIC POSTRHEUMATIC ARTHROPATHY, UNSPECIFIED KNEE
C4270415|T046|T83.728A|ICD10CM|EXPOSURE OF OTHER IMPLANTED MESH INTO ORGAN OR TISSUE, INITIAL ENCOUNTER|EXPOSURE OF OTHER IMPLANTED MESH INTO ORGAN OR TISSUE, INIT
C2832319|T037|S06.363S|ICD10CM|TRAUMATIC HEMORRHAGE OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF 1 HOURS TO 5 HOURS 59 MINUTES, SEQUELA|TRAUM HEMOR CEREB, W LOC OF 1-5 HRS 59 MINUTES, SEQUELA
C2886735|T037|T79.5XXA|ICD10CM|TRAUMATIC ANURIA, INITIAL ENCOUNTER|TRAUMATIC ANURIA, INITIAL ENCOUNTER
C2875155|T047|G43.401|ICD10CM|HEMIPLEGIC MIGRAINE, NOT INTRACTABLE, WITH STATUS MIGRAINOSUS|HEMIPLEGIC MIGRAINE, NOT INTRACTABLE, W STATUS MIGRAINOSUS
C2895323|T037|M48.53XA|ICD10CM|COLLAPSED VERTEBRA, NOT ELSEWHERE CLASSIFIED, CERVICOTHORACIC REGION, INITIAL ENCOUNTER FOR FRACTURE|COLLAPSED VERTEBRA, NEC, CERVICOTHORACIC REGION, INIT
C2875156|T047|G43.409|ICD10CM|HEMIPLEGIC MIGRAINE, NOT INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|HEMIPLEGIC MIGRAINE, NOT INTRACTABLE, W/O STATUS MIGRAINOSUS
C0751560|T191|C09.9|DMDICD10|MALIGNANT NEOPLASM OF TONSIL, UNSPECIFIED|BOESARTIGE NEUBILDUNG: TONSILLE, NICHT NAEHER BEZEICHNET
C2874641|T048|F15.19|ICD10CM|OTHER STIMULANT ABUSE WITH UNSPECIFIED STIMULANT-INDUCED DISORDER|OTHER STIMULANT ABUSE WITH UNSP STIMULANT-INDUCED DISORDER
C4268246|T048|F15.14|ICD10CM|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED MOOD DISORDER|AMPHETAMINE OR OTHER STIMULANT USE DISORDER, MILD, WITH AMPHETAMINE OR OTHER STIMULANT INDUCED DEPRESSIVE DISORDER
C4065855|T048||ICD10CM|CONVERSION DISORDER WITH SENSORY SYMPTOM OR DEFICIT
C2874952|T048|F44.7|ICD10CM|CONVERSION DISORDER WITH MIXED SYMPTOM PRESENTATION|CONVERSION DISORDER WITH MIXED SYMPTOM PRESENTATION
C4509115|T048|F44.4|ICD10CM|CONVERSION DISORDER WITH MOTOR SYMPTOM OR DEFICIT|CONVERSION DISORDER WITH WEAKNESS/PARALYSIS
C4065854|T048||ICD10CM|CONVERSION DISORDER WITH SEIZURES OR CONVULSIONS
C0349449|T048|F44.2|DMDICD10|DISSOCIATIVE STUPOR|DISSOZIATIVER STUPOR
C0236795|T048|F44.0|DMDICD10|DISSOCIATIVE AMNESIA|DISSOZIATIVE AMNESIE
C4237105|T048|F44.1|ICD10CM|DISSOCIATIVE FUGUE|DISSOCIATIVE AMNESIA WITH DISSOCIATIVE FUGUE
C2835768|T037|S24.104A|ICD10CM|UNSPECIFIED INJURY AT T11-T12 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY AT T11-T12 LEVEL OF THORACIC SPINAL CORD, INIT
C2876870|T037|T37.3X2S|ICD10CM|POISONING BY OTHER ANTIPROTOZOAL DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH ANTIPROTOZOAL DRUGS, SELF-HARM, SEQUELA
C2835857|T037|S24.159A|ICD10CM|OTHER INCOMPLETE LESION AT UNSPECIFIED LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|OTH INCMPL LESION AT UNSP LEVEL OF THOR SPINAL CORD, INIT
C2835769|T037|S24.104D|ICD10CM|UNSPECIFIED INJURY AT T11-T12 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY AT T11-T12 LEVEL OF THORACIC SPINAL CORD, SUBS
C1442976|T048|F44|DMDICD10|DISSOCIATIVE AND CONVERSION DISORDER, UNSPECIFIED|DISSOZIATIVE STOERUNGEN [KONVERSIONSSTOERUNGEN]
C2900579|T047|M81.0|ICD10CM|AGE-RELATED OSTEOPOROSIS WITHOUT CURRENT PATHOLOGICAL FRACTURE|AGE-RELATED OSTEOPOROSIS W/O CURRENT PATHOLOGICAL FRACTURE
C0451868|T047|M81.6|DMDICD10|LOCALIZED OSTEOPOROSIS [LEQUESNE]|LOKALISIERTE OSTEOPOROSE [LEQUESNE]
C2900586|T046|M81.8|ICD10CM|OTHER OSTEOPOROSIS WITHOUT CURRENT PATHOLOGICAL FRACTURE|OTHER OSTEOPOROSIS WITHOUT CURRENT PATHOLOGICAL FRACTURE
C2835770|T037|S24.104S|ICD10CM|UNSPECIFIED INJURY AT T11-T12 LEVEL OF THORACIC SPINAL CORD, SEQUELA|UNSP INJURY AT T11-T12, SEQUELA
C2833928|T037|S14.123D|ICD10CM|CENTRAL CORD SYNDROME AT C3 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|CENTRAL CORD SYNDROME AT C3, SUBS
C2845961|T191|C78.7|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF LIVER AND INTRAHEPATIC BILE DUCT|SECONDARY MALIG NEOPLASM OF LIVER AND INTRAHEPATIC BILE DUCT
C2883938|T037|T50.Z12A|ICD10CM|POISONING BY IMMUNOGLOBULIN, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY IMMUNOGLOBULIN, INTENTIONAL SELF-HARM, INIT
C4269328|T037|S02.11HA|ICD10CM|OTHER FRACTURE OF OCCIPUT, LEFT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTHER FRACTURE OF OCCIPUT, LEFT SIDE, INIT
C4269329|T037|S02.11HB|ICD10CM|OTHER FRACTURE OF OCCIPUT, LEFT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTHER FRACTURE OF OCCIPUT, LEFT SIDE, 7THB
C0477969|T019|Q01.8|DMDICD10|ENCEPHALOCELE OF OTHER SITES|ENZEPHALOZELE SONSTIGER LOKALISATIONEN
C2854085|T191|C90.32|ICD10CM|SOLITARY PLASMACYTOMA IN RELAPSE|SOLITARY PLASMACYTOMA IN RELAPSE
C4269333|T037|S02.11HS|ICD10CM|OTHER FRACTURE OF OCCIPUT, LEFT SIDE, SEQUELA|OTHER FRACTURE OF OCCIPUT, LEFT SIDE, SEQUELA
C0431289|T019|Q01.0|DMDICD10|FRONTAL ENCEPHALOCELE|FRONTALE ENZEPHALOZELE
C0431291|T019|Q01.1|DMDICD10|NASOFRONTAL ENCEPHALOCELE|NASOFRONTALE ENZEPHALOZELE
C0014067|T019|Q01.2|DMDICD10|OCCIPITAL ENCEPHALOCELE|OKZIPITALE ENZEPHALOZELE
C2857395|T037|S72.133B|ICD10CM|DISPLACED APOPHYSEAL FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPLACED APOPHYSEAL FX UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2857396|T037|S72.133C|ICD10CM|DISPLACED APOPHYSEAL FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL APOPHYSEAL FX UNSP FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2857394|T037|S72.133A|ICD10CM|DISPLACED APOPHYSEAL FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED APOPHYSEAL FRACTURE OF UNSP FEMUR, INIT
C2838705|T037|S34.139S|ICD10CM|UNSPECIFIED INJURY TO SACRAL SPINAL CORD, SEQUELA|UNSPECIFIED INJURY TO SACRAL SPINAL CORD, SEQUELA
C2889177|T047|M05.239|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF UNSP WRIST
C2882763|T047|I70.329|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, UNSPECIFIED EXTREMITY|ATHSCL UNSP TYPE BYPASS OF THE EXTRM W REST PAIN, UNSP EXTRM
C2882762|T047|I70.328|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, OTHER EXTREMITY|ATHSCL UNSP TYPE BYPASS OF THE EXTRM W REST PAIN, OTH EXTRM
C2882761|T047|I70.323|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, BILATERAL LEGS|ATHSCL UNSP TYPE BYPASS OF THE EXTRM W REST PAIN, BI LEGS
C2882760|T047|I70.322|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, LEFT LEG|ATHSCL UNSP TYPE BYPASS OF THE EXTRM W REST PAIN, LEFT LEG
C2882759|T047|I70.321|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, RIGHT LEG|ATHSCL UNSP TYPE BYPASS OF THE EXTRM W REST PAIN, RIGHT LEG
C2889176|T047|M05.232|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT WRIST|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF LEFT WRIST
C2869874|T037|S98.321A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT MIDFOOT, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF RIGHT MIDFOOT, INIT ENCNTR
C2869876|T037|S98.321S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT MIDFOOT, SEQUELA|PARTIAL TRAUMATIC AMPUTATION OF RIGHT MIDFOOT, SEQUELA
C2876234|T037|T32.98|ICD10CM|CORROSIONS INVOLVING 90% OR MORE OF BODY SURFACE WITH 80-89% THIRD DEGREE CORROSION|CORROS 90%/MORE OF BODY SURFACE W 80-89% THIRD DEGREE CORROS
C2837640|T037|S32.052B|ICD10CM|UNSTABLE BURST FRACTURE OF FIFTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSTABLE BURST FX FIFTH LUM VERTEBRA, INIT FOR OPN FX
C2833466|T037|S12.430B|ICD10CM|UNSPECIFIED TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP TRAUM DISPL SPONDYLOLYSIS OF 5TH CERVCAL VERT, 7THB
C2885594|T037|T63.392S|ICD10CM|TOXIC EFFECT OF VENOM OF OTHER SPIDER, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF SPIDER, SELF-HARM, SEQUELA
C4269249|T037|S02.109S|ICD10CM|FRACTURE OF BASE OF SKULL, UNSPECIFIED SIDE, SEQUELA|FRACTURE OF BASE OF SKULL, UNSPECIFIED SIDE, SEQUELA
C2890203|T037|T83.010A|ICD10CM|BREAKDOWN (MECHANICAL) OF CYSTOSTOMY CATHETER, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF CYSTOSTOMY CATHETER, INIT ENCNTR
C2885592|T037|T63.392A|ICD10CM|TOXIC EFFECT OF VENOM OF OTHER SPIDER, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF SPIDER, INTENTIONAL SELF-HARM, INIT
C2902741|T037|M96.671|ICD10CM|FRACTURE OF TIBIA OR FIBULA FOLLOWING INSERTION OF ORTHOPEDIC IMPLANT, JOINT PROSTHESIS, OR BONE PLATE, RIGHT LEG|FX TIB/FIB FOL INSRT ORTHO IMPLNT/PROSTH/BONE PLT, RIGHT LEG
C2902742|T037|M96.672|ICD10CM|FRACTURE OF TIBIA OR FIBULA FOLLOWING INSERTION OF ORTHOPEDIC IMPLANT, JOINT PROSTHESIS, OR BONE PLATE, LEFT LEG|FX TIB/FIB FOL INSRT ORTHO IMPLNT/PROSTH/BONE PLT, LEFT LEG
C2835413|T037|S22.071A|ICD10CM|STABLE BURST FRACTURE OF T9-T10 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|STABLE BURST FRACTURE OF T9-T10 VERTEBRA, INIT FOR CLOS FX
C2835414|T037|S22.071B|ICD10CM|STABLE BURST FRACTURE OF T9-T10 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|STABLE BURST FRACTURE OF T9-T10 VERTEBRA, INIT FOR OPN FX
C2902743|T037|M96.679|ICD10CM|FRACTURE OF TIBIA OR FIBULA FOLLOWING INSERTION OF ORTHOPEDIC IMPLANT, JOINT PROSTHESIS, OR BONE PLATE, UNSPECIFIED LEG|FX TIB/FIB FOL INSRT ORTHO IMPLNT/PROSTH/BONE PLT, UNSP LEG
C4269244|T037|S02.109A|ICD10CM|FRACTURE OF BASE OF SKULL, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF BASE OF SKULL, UNSPECIFIED SIDE, INIT
C2832643|T037|S06.893A|ICD10CM|OTHER SPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|INTCRAN INJ W LOSS OF CONSCIOUSNESS OF 1-5 HRS 59 MIN, INIT
C2901938|T046|M87.012|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF LEFT SHOULDER|IDIOPATHIC ASEPTIC NECROSIS OF LEFT SHOULDER
C4509298|T047|L97.318|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT ANKLE WITH OTHER SPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF RIGHT ANKLE WITH OTH SEVERITY
C2888687|T047|L97.319|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT ANKLE WITH UNSPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF RIGHT ANKLE WITH UNSP SEVERITY
C4509297|T047|L97.316|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT ANKLE WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULCER OF R ANKLE WITH BONE INVL W/O EVD OF NECR
C2888686|T047|L97.314|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT ANKLE WITH NECROSIS OF BONE|NON-PRESSURE CHRONIC ULCER OF RIGHT ANKLE W NECROSIS OF BONE
C4509296|T047|L97.315|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT ANKLE WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULCER OF R ANKLE WITH MSL INVL W/O EVD OF NECR
C2888684|T047|L97.312|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT ANKLE WITH FAT LAYER EXPOSED|NON-PRS CHRONIC ULCER OF RIGHT ANKLE W FAT LAYER EXPOSED
C2888685|T047|L97.313|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT ANKLE WITH NECROSIS OF MUSCLE|NON-PRS CHRONIC ULCER OF RIGHT ANKLE W NECROSIS OF MUSCLE
C2901939|T046|M87.019|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED SHOULDER|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED SHOULDER
C2888683|T047|L97.311|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT ANKLE LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHRONIC ULCER OF RIGHT ANKLE LIMITED TO BRKDWN SKIN
C2869808|T037|S98.131D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF ONE RIGHT LESSER TOE, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF ONE RIGHT LESSER TOE, SUBS
C2832525|T037|S06.6X4A|ICD10CM|TRAUMATIC SUBARACHNOID HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|TRAUM SUBRAC HEM W LOC OF 6 HOURS TO 24 HOURS, INIT
C2883082|T047|I82.210|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF SUPERIOR VENA CAVA|ACUTE EMBOLISM AND THROMBOSIS OF SUPERIOR VENA CAVA
C2883083|T047|I82.211|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF SUPERIOR VENA CAVA|CHRONIC EMBOLISM AND THROMBOSIS OF SUPERIOR VENA CAVA
C2890354|T037|T83.490A|ICD10CM|OTHER MECHANICAL COMPLICATION OF IMPLANTED PENILE PROSTHESIS, INITIAL ENCOUNTER|MECH COMPL OF IMPLANTED PENILE PROSTHESIS, INITIAL ENCOUNTER
C2838450|T037|S32.614A|ICD10CM|NONDISPLACED AVULSION FRACTURE OF RIGHT ISCHIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED AVULSION FRACTURE OF RIGHT ISCHIUM, INIT
C2838451|T037|S32.614B|ICD10CM|NONDISPLACED AVULSION FRACTURE OF RIGHT ISCHIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP AVULSION FRACTURE OF RIGHT ISCHIUM, INIT FOR OPN FX
C2837861|T037|S32.316B|ICD10CM|NONDISPLACED AVULSION FRACTURE OF UNSPECIFIED ILIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP AVULSION FRACTURE OF UNSP ILIUM, INIT FOR OPN FX
C2860050|T037|S79.001A|ICD10CM|UNSPECIFIED PHYSEAL FRACTURE OF UPPER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP PHYSEAL FRACTURE OF UPPER END OF RIGHT FEMUR, INIT
C0271847|T047|N25.81|ICD10CM|SECONDARY HYPERPARATHYROIDISM OF RENAL ORIGIN|SECONDARY HYPERPARATHYROIDISM OF RENAL ORIGIN
C4267917|T047|E08.3491|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|DIABETES WITH SEVERE NONP RTNOP WITHOUT MACULAR EDEMA, R EYE
C2856073|T037|S68.627S|ICD10CM|PARTIAL TRAUMATIC TRANSPHALANGEAL AMPUTATION OF LEFT LITTLE FINGER, SEQUELA|PARTIAL TRAUMATIC TRNSPHAL AMP OF L LITTLE FINGER, SEQUELA
C2838496|T037|S32.810B|ICD10CM|MULTIPLE FRACTURES OF PELVIS WITH STABLE DISRUPTION OF PELVIC RING, INITIAL ENCOUNTER FOR OPEN FRACTURE|MULT FX OF PELV W STABLE DISRUPT OF PELV RING, 7THB
C2896662|T046|M80.811A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, RIGHT SHOULDER, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, R SHOULDER, INIT
C2858954|T037|S72.471A|ICD10CM|TORUS FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TORUS FRACTURE OF LOWER END OF RIGHT FEMUR, INIT FOR CLOS FX
C2834062|T037|S14.158S|ICD10CM|OTHER INCOMPLETE LESION AT C8 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|OTH INCOMPLETE LESION AT C8, SEQUELA
C2845973|T191|C79.72|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF LEFT ADRENAL GLAND|SECONDARY MALIGNANT NEOPLASM OF LEFT ADRENAL GLAND
C2845972|T191|C79.71|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF RIGHT ADRENAL GLAND|SECONDARY MALIGNANT NEOPLASM OF RIGHT ADRENAL GLAND
C2845971|T191|C79.70|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF UNSPECIFIED ADRENAL GLAND|SECONDARY MALIGNANT NEOPLASM OF UNSPECIFIED ADRENAL GLAND
C2834061|T037|S14.158D|ICD10CM|OTHER INCOMPLETE LESION AT C8 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|OTH INCOMPLETE LESION AT C8, SUBS
C2878611|T037|T43.622A|ICD10CM|POISONING BY AMPHETAMINES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY AMPHETAMINES, INTENTIONAL SELF-HARM, INIT
C2834060|T037|S14.158A|ICD10CM|OTHER INCOMPLETE LESION AT C8 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|OTH INCOMPLETE LESION AT C8, INIT
C0343453|T047|A26.7|DMDICD10|ERYSIPELOTHRIX SEPSIS|ERYSIPELOTHRIX-SEPSIS
C2858938|T037|S72.466C|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP SUPRCNDL FX W INTRCNDL EXTN LOW END UNSP FEMR, 7THC
C2891336|T047||ICD10CM|NECROSIS OF AMPUTATION STUMP, LEFT UPPER EXTREMITY
C2879259|T037|T45.622S|ICD10CM|POISONING BY HEMOSTATIC DRUG, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY HEMOSTATIC DRUG, INTENTIONAL SELF-HARM, SEQUELA
C2860222|T037|S79.149A|ICD10CM|SALTER-HARRIS TYPE IV PHYSEAL FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SLTR-HARIS TYPE IV PHYSEAL FX LOWER END OF UNSP FEMUR, INIT
C2884004|T037|T51.1X2S|ICD10CM|TOXIC EFFECT OF METHANOL, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF METHANOL, INTENTIONAL SELF-HARM, SEQUELA
C0477402|T047|G61|DMDICD10|INFLAMMATORY POLYNEUROPATHY, UNSPECIFIED|POLYNEURITIS
C2884849|T037|T59.1X2A|ICD10CM|TOXIC EFFECT OF SULFUR DIOXIDE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF SULFUR DIOXIDE, INTENTIONAL SELF-HARM, INIT
C2876227|T037|T32.91|ICD10CM|CORROSIONS INVOLVING 90% OR MORE OF BODY SURFACE WITH 10-19% THIRD DEGREE CORROSION|CORROS 90%/MORE OF BODY SURFACE W 10-19% THIRD DEGREE CORROS
C2902738|T037|M96.662|ICD10CM|FRACTURE OF FEMUR FOLLOWING INSERTION OF ORTHOPEDIC IMPLANT, JOINT PROSTHESIS, OR BONE PLATE, LEFT LEG|FX FEMUR FOL INSRT ORTHO IMPLNT/PROSTH/BONE PLT, LEFT LEG
C2875304|T047|G61.0|ICD10CM|GUILLAIN-BARRE SYNDROME|ACUTE (POST-)INFECTIVE POLYNEURITIS
C0451648|T047|G61.1|DMDICD10|SERUM NEUROPATHY|SERUMPOLYNEUROPATHIE
C2837721|T037|S32.129B|ICD10CM|UNSPECIFIED ZONE II FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP ZONE II FRACTURE OF SACRUM, INIT FOR OPN FX
C2902737|T037|M96.661|ICD10CM|FRACTURE OF FEMUR FOLLOWING INSERTION OF ORTHOPEDIC IMPLANT, JOINT PROSTHESIS, OR BONE PLATE, RIGHT LEG|FX FEMUR FOL INSRT ORTHO IMPLNT/PROSTH/BONE PLT, RIGHT LEG
C0155858|T047|J15.8|DMDICD10|PNEUMONIA DUE TO OTHER SPECIFIED BACTERIA|SONSTIGE BAKTERIELLE PNEUMONIE
C0375326|T047|J15.4|DMDICD10|PNEUMONIA DUE TO OTHER STREPTOCOCCI|PNEUMONIE DURCH SONSTIGE STREPTOKOKKEN
C0276089|T047|J15.5|DMDICD10|PNEUMONIA DUE TO ESCHERICHIA COLI|PNEUMONIE DURCH ESCHERICHIA COLI
C0865782|T047|J15.6|ICD10CM|PNEUMONIA DUE TO OTHER GRAM-NEGATIVE BACTERIA|PNEUMONIA DUE TO SERRATIA MARCESCENS
C2879593|T037|T46.8X2A|ICD10CM|POISONING BY ANTIVARICOSE DRUGS, INCLUDING SCLEROSING AGENTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY ANTIVARIC DRUGS, INC SCLER AGENTS, SELF-HARM, INIT
C0519030|T047|B96.1|DMDICD10|PNEUMONIA DUE TO KLEBSIELLA PNEUMONIAE|KLEBSIELLA PNEUMONIAE [K. PNEUMONIAE] ALS URSACHE VON KRANKHEITEN, DIE IN ANDEREN KAPITELN KLASSIFIZIERT SIND
C0155860|T047|J15.1|DMDICD10|PNEUMONIA DUE TO PSEUDOMONAS|PNEUMONIE DURCH PSEUDOMONAS
C0348801|T047|J15.3|DMDICD10|PNEUMONIA DUE TO STREPTOCOCCUS, GROUP B|PNEUMONIE DURCH STREPTOKOKKEN DER GRUPPE B
C2879646|T037|T46.992S|ICD10CM|POISONING BY OTHER AGENTS PRIMARILY AFFECTING THE CARDIOVASCULAR SYSTEM, INTENTIONAL SELF-HARM, SEQUELA|POISN BY OTH AGENTS AFF THE CARDIOVASC SYS, SLF-HRM, SEQUELA
C0856761|T047|I82.0|DMDICD10|BUDD-CHIARI SYNDROME|BUDD-CHIARI-SYNDROM
C0155776|T046|I82.3|DMDICD10|EMBOLISM AND THROMBOSIS OF RENAL VEIN|EMBOLIE UND THROMBOSE DER NIERENVENE
C2878613|T037|T43.622S|ICD10CM|POISONING BY AMPHETAMINES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY AMPHETAMINES, INTENTIONAL SELF-HARM, SEQUELA
C2890429|T037|T84.020A|ICD10CM|DISLOCATION OF INTERNAL RIGHT HIP PROSTHESIS, INITIAL ENCOUNTER|DISLOCATION OF INTERNAL RIGHT HIP PROSTHESIS, INIT ENCNTR
C2884833|T037|T59.0X2A|ICD10CM|TOXIC EFFECT OF NITROGEN OXIDES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF NITROGEN OXIDES, INTENTIONAL SELF-HARM, INIT
C0221046|T047|G90.01|ICD10CM|CAROTID SINUS SYNCOPE|CAROTID SINUS SYNDROME
C2876229|T037|T32.93|ICD10CM|CORROSIONS INVOLVING 90% OR MORE OF BODY SURFACE WITH 30-39% THIRD DEGREE CORROSION|CORROS 90%/MORE OF BODY SURFACE W 30-39% THIRD DEGREE CORROS
C2349411|T047|G90.09|ICD10CM|OTHER IDIOPATHIC PERIPHERAL AUTONOMIC NEUROPATHY|OTHER IDIOPATHIC PERIPHERAL AUTONOMIC NEUROPATHY
C2838655|T037|S34.114S|ICD10CM|COMPLETE LESION OF L4 LEVEL OF LUMBAR SPINAL CORD, SEQUELA|COMPLETE LESION OF L4 LEVEL OF LUMBAR SPINAL CORD, SEQUELA
C2869871|T037|S98.319S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED MIDFOOT, SEQUELA|COMPLETE TRAUMATIC AMPUTATION OF UNSP MIDFOOT, SEQUELA
C2875115|T047|G40.411|ICD10CM|OTHER GENERALIZED EPILEPSY AND EPILEPTIC SYNDROMES, INTRACTABLE, WITH STATUS EPILEPTICUS|OTH GENERALIZED EPILEPSY, INTRACTABLE, W STATUS EPILEPTICUS
C2874784|T048|F18.980|ICD10CM|INHALANT USE, UNSPECIFIED WITH INHALANT-INDUCED ANXIETY DISORDER|INHALANT USE, UNSP WITH INHALANT-INDUCED ANXIETY DISORDER
C2859977|T037|S78.012S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEFT HIP JOINT, SEQUELA|COMPLETE TRAUMATIC AMPUTATION AT LEFT HIP JOINT, SEQUELA
C2896626|T046|M80.072A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, LEFT ANKLE AND FOOT, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, LEFT ANK/FT, INIT
C4237514|T048|F18.988|ICD10CM|INHALANT USE, UNSPECIFIED WITH OTHER INHALANT-INDUCED DISORDER|INHALANT-INDUCED MILD NEUROCOGNITIVE DISORDER
C2859976|T037|S78.012D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEFT HIP JOINT, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION AT LEFT HIP JOINT, SUBS ENCNTR
C0242670|T047||ICD10CM|PERSISTENT VEGETATIVE STATE
C2859975|T037|S78.012A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEFT HIP JOINT, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION AT LEFT HIP JOINT, INIT ENCNTR
C2838129|T037|S32.436B|ICD10CM|NONDISPLACED FRACTURE OF ANTERIOR COLUMN [ILIOPUBIC] OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP FX OF ANT COLUMN OF UNSP ACETAB, INIT FOR OPN FX
C2838128|T037|S32.436A|ICD10CM|NONDISPLACED FRACTURE OF ANTERIOR COLUMN [ILIOPUBIC] OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF ANTERIOR COLUMN OF UNSP ACETABULUM, INIT
C2838308|T037|S32.481A|ICD10CM|DISPLACED DOME FRACTURE OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED DOME FRACTURE OF RIGHT ACETABULUM, INIT
C2838309|T037|S32.481B|ICD10CM|DISPLACED DOME FRACTURE OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISPLACED DOME FRACTURE OF RIGHT ACETABULUM, INIT FOR OPN FX
C2832690|T037|S06.9X4S|ICD10CM|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|UNSP INTRACRANIAL INJURY W LOC OF 6-24 HRS, SEQUELA
C2884851|T037|T59.1X2S|ICD10CM|TOXIC EFFECT OF SULFUR DIOXIDE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF SULFUR DIOXIDE, SELF-HARM, SEQUELA
C4267913|T047|E08.3411|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|DIABETES WITH SEVERE NONP RTNOP WITH MACULAR EDEMA, R EYE
C4267914|T047|E08.3412|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|DIABETES WITH SEVERE NONP RTNOP WITH MACULAR EDEMA, LEFT EYE
C4267915|T047|E08.3413|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|DIABETES WITH SEVERE NONP RTNOP WITH MACULAR EDEMA, BI
C2879749|T037|T47.3X2S|ICD10CM|POISONING BY SALINE AND OSMOTIC LAXATIVES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY SALINE AND OSMOTIC LAXTV, SELF-HARM, SEQUELA
C2882961|T047|I70.662|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, LEFT LEG|ATHSCL NONBIOL BYPASS OF THE EXTRM W GANGRENE, LEFT LEG
C2887312|T047|I87.333|ICD10CM|CHRONIC VENOUS HYPERTENSION (IDIOPATHIC) WITH ULCER AND INFLAMMATION OF BILATERAL LOWER EXTREMITY|CHRONIC VENOUS HTN W ULCER AND INFLAM OF BILATERAL LOW EXTRM
C2887310|T047|I87.331|ICD10CM|CHRONIC VENOUS HYPERTENSION (IDIOPATHIC) WITH ULCER AND INFLAMMATION OF RIGHT LOWER EXTREMITY|CHRONIC VENOUS HTN W ULCER AND INFLAMMATION OF R LOW EXTREM
C2832688|T037|S06.9X4A|ICD10CM|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|UNSP INTRACRANIAL INJURY W LOC OF 6 HOURS TO 24 HOURS, INIT
C2905743|T037|X77.8XXD|ICD10CM|INTENTIONAL SELF-HARM BY OTHER HOT OBJECTS, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY OTHER HOT OBJECTS, SUBS ENCNTR
C2854031|T191|C85.18|ICD10CM|UNSPECIFIED B-CELL LYMPHOMA, LYMPH NODES OF MULTIPLE SITES|UNSPECIFIED B-CELL LYMPHOMA, LYMPH NODES OF MULTIPLE SITES
C2854032|T191|C85.19|ICD10CM|UNSPECIFIED B-CELL LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES|UNSP B-CELL LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES
C2854027|T191|C85.14|ICD10CM|UNSPECIFIED B-CELL LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB|UNSP B-CELL LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB
C2854028|T191|C85.15|ICD10CM|UNSPECIFIED B-CELL LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|UNSP B-CELL LYMPHOMA, NODES OF ING REGION AND LOWER LIMB
C2854029|T191|C85.16|ICD10CM|UNSPECIFIED B-CELL LYMPHOMA, INTRAPELVIC LYMPH NODES|UNSPECIFIED B-CELL LYMPHOMA, INTRAPELVIC LYMPH NODES
C2854030|T191|C85.17|ICD10CM|UNSPECIFIED B-CELL LYMPHOMA, SPLEEN|UNSPECIFIED B-CELL LYMPHOMA, SPLEEN
C2854023|T191|C85.10|ICD10CM|UNSPECIFIED B-CELL LYMPHOMA, UNSPECIFIED SITE|UNSPECIFIED B-CELL LYMPHOMA, UNSPECIFIED SITE
C2854024|T191|C85.11|ICD10CM|UNSPECIFIED B-CELL LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK|UNSP B-CELL LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK
C2854025|T191|C85.12|ICD10CM|UNSPECIFIED B-CELL LYMPHOMA, INTRATHORACIC LYMPH NODES|UNSPECIFIED B-CELL LYMPHOMA, INTRATHORACIC LYMPH NODES
C2854026|T191|C85.13|ICD10CM|UNSPECIFIED B-CELL LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES|UNSPECIFIED B-CELL LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES
C2888854|T047|M00.171|ICD10CM|PNEUMOCOCCAL ARTHRITIS, RIGHT ANKLE AND FOOT|PNEUMOCOCCAL ARTHRITIS, RIGHT ANKLE AND FOOT
C2888855|T047|M00.172|ICD10CM|PNEUMOCOCCAL ARTHRITIS, LEFT ANKLE AND FOOT|PNEUMOCOCCAL ARTHRITIS, LEFT ANKLE AND FOOT
C4268277|T048|F18.188|ICD10CM|INHALANT ABUSE WITH OTHER INHALANT-INDUCED DISORDER|INHALANT USE DISORDER, MILD, WITH INHALANT INDUCED MILD NEUROCOGNITIVE DISORDER
C2890801|T037|T84.50XA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO UNSPECIFIED INTERNAL JOINT PROSTHESIS, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO UNSP INT JOINT PROSTH, INIT
C2888856|T047|M00.179|ICD10CM|PNEUMOCOCCAL ARTHRITIS, UNSPECIFIED ANKLE AND FOOT|PNEUMOCOCCAL ARTHRITIS, UNSPECIFIED ANKLE AND FOOT
C2874756|T048|F18.180|ICD10CM|INHALANT ABUSE WITH INHALANT-INDUCED ANXIETY DISORDER|INHALANT ABUSE WITH INHALANT-INDUCED ANXIETY DISORDER
C2891163|T037|T85.621S|ICD10CM|DISPLACEMENT OF INTRAPERITONEAL DIALYSIS CATHETER, SEQUELA|DISPLACEMENT OF INTRAPERITONEAL DIALYSIS CATHETER, SEQUELA
C2890817|T037|T84.54XA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL LEFT KNEE PROSTHESIS, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INTERNAL LEFT KNEE PROSTH, INIT
C2886762|T037|T79.A21A|ICD10CM|TRAUMATIC COMPARTMENT SYNDROME OF RIGHT LOWER EXTREMITY, INITIAL ENCOUNTER|TRAUMATIC COMPARTMENT SYNDROME OF R LOW EXTREM, INIT
C2891162|T037|T85.621D|ICD10CM|DISPLACEMENT OF INTRAPERITONEAL DIALYSIS CATHETER, SUBSEQUENT ENCOUNTER|DISPLACEMENT OF INTRAPERITONEAL DIALYSIS CATHETER, SUBS
C2891161|T037|T85.621A|ICD10CM|DISPLACEMENT OF INTRAPERITONEAL DIALYSIS CATHETER, INITIAL ENCOUNTER|DISPLACEMENT OF INTRAPERITONEAL DIALYSIS CATHETER, INIT
C3263978|T047|G40.811|ICD10CM|LENNOX-GASTAUT SYNDROME, NOT INTRACTABLE, WITH STATUS EPILEPTICUS|LENNOX-GASTAUT SYNDROME, NOT INTRACTABLE, W STAT EPI
C3263979|T047|G40.812|ICD10CM|LENNOX-GASTAUT SYNDROME, NOT INTRACTABLE, WITHOUT STATUS EPILEPTICUS|LENNOX-GASTAUT SYNDROME, NOT INTRACTABLE, W/O STAT EPI
C3263980|T047|G40.813|ICD10CM|LENNOX-GASTAUT SYNDROME, INTRACTABLE, WITH STATUS EPILEPTICUS|LENNOX-GASTAUT SYNDROME, INTRACTABLE, W STATUS EPILEPTICUS
C3263981|T047|G40.814|ICD10CM|LENNOX-GASTAUT SYNDROME, INTRACTABLE, WITHOUT STATUS EPILEPTICUS|LENNOX-GASTAUT SYNDROME, INTRACTABLE, W/O STATUS EPILEPTICUS
C2905720|T037|X75.XXXD|ICD10CM|INTENTIONAL SELF-HARM BY EXPLOSIVE MATERIAL, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY EXPLOSIVE MATERIAL, SUBS ENCNTR
C2905719|T037|X75.XXXA|ICD10CM|INTENTIONAL SELF-HARM BY EXPLOSIVE MATERIAL, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY EXPLOSIVE MATERIAL, INIT ENCNTR
C2856587|T037|S72.021B|ICD10CM|DISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF EPIPHY (SEPARATION) (UPPER) OF R FEMR, 7THB
C2855993|T037|S68.522S|ICD10CM|PARTIAL TRAUMATIC TRANSPHALANGEAL AMPUTATION OF LEFT THUMB, SEQUELA|PARTIAL TRAUMATIC TRNSPHAL AMPUTATION OF LEFT THUMB, SEQUELA
C2856586|T037|S72.021A|ICD10CM|DISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF EPIPHYSIS (SEPARATION) (UPPER) OF R FEMUR, INIT
C2873766|T047||ICD10CM|SICKLE-CELL THALASSEMIA WITH ACUTE CHEST SYNDROME
C2873767|T047||ICD10CM|SICKLE-CELL THALASSEMIA WITH SPLENIC SEQUESTRATION
C1260395|T047|D57.419|ICD10CM|SICKLE-CELL THALASSEMIA WITH CRISIS, UNSPECIFIED|SICKLE-CELL THALASSEMIA WITH CRISIS, UNSPECIFIED
C2857498|T037|S72.143C|ICD10CM|DISPLACED INTERTROCHANTERIC FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL INTERTROCH FX UNSP FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2857497|T037|S72.143B|ICD10CM|DISPLACED INTERTROCHANTERIC FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPLACED INTERTROCH FX UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2901851|T047|M86.339|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, UNSPECIFIED RADIUS AND ULNA|CHRONIC MULTIFOCAL OSTEOMYELITIS, UNSP RADIUS AND ULNA
C2833908|T037|S14.117S|ICD10CM|COMPLETE LESION AT C7 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|COMPLETE LESION AT C7 LEVEL OF CERVICAL SPINAL CORD, SEQUELA
C0024523|T047|K90.9|DMDICD10|INTESTINAL MALABSORPTION, UNSPECIFIED|INTESTINALE MALABSORPTION, NICHT NAEHER BEZEICHNET
C2901849|T047|M86.331|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, RIGHT RADIUS AND ULNA|CHRONIC MULTIFOCAL OSTEOMYELITIS, RIGHT RADIUS AND ULNA
C2885524|T037|T63.302A|ICD10CM|TOXIC EFFECT OF UNSPECIFIED SPIDER VENOM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF UNSP SPIDER VENOM, SELF-HARM, INIT
C2901850|T047|M86.332|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, LEFT RADIUS AND ULNA|CHRONIC MULTIFOCAL OSTEOMYELITIS, LEFT RADIUS AND ULNA
C4509268|T047|K90.0|ICD10CM|CELIAC DISEASE|CELIAC GLUTEN-SENSITIVE ENTEROPATHY
C0205707|T047||ICD10CM|TROPICAL SPRUE
C0494805|T047|K90.2|DMDICD10|BLIND LOOP SYNDROME, NOT ELSEWHERE CLASSIFIED|SYNDROM DER BLINDEN SCHLINGE, ANDERENORTS NICHT KLASSIFIZIERT
C0152166|T047|K90.3|DMDICD10|PANCREATIC STEATORRHEA|PANKREATOGENE STEATORRHOE
C2832144|T037|S06.322A|ICD10CM|CONTUSION AND LACERATION OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|CONTUS/LAC LEFT CEREBRUM W LOC OF 31-59 MIN, INIT
C2855980|T037|S68.512S|ICD10CM|COMPLETE TRAUMATIC TRANSPHALANGEAL AMPUTATION OF LEFT THUMB, SEQUELA|COMPLETE TRAUMATIC TRNSPHAL AMP OF LEFT THUMB, SEQUELA
C2874051|T047|E10.51|ICD10CM|TYPE 1 DIABETES MELLITUS WITH DIABETIC PERIPHERAL ANGIOPATHY WITHOUT GANGRENE|TYPE 1 DIABETES W DIABETIC PERIPHERAL ANGIOPATH W/O GANGRENE
C2874053|T047|E10.52|ICD10CM|TYPE 1 DIABETES MELLITUS WITH DIABETIC PERIPHERAL ANGIOPATHY WITH GANGRENE|TYPE 1 DIABETES W DIABETIC PERIPHERAL ANGIOPATHY W GANGRENE
C0432452|T047|Q95.2|DMDICD10|BALANCED AUTOSOMAL REARRANGEMENT IN ABNORMAL INDIVIDUAL|BALANCIERTES REARRANGEMENT DER AUTOSOMEN BEIM ABNORMEN INDIVIDUUM
C2874054|T047|E10.59|ICD10CM|TYPE 1 DIABETES MELLITUS WITH OTHER CIRCULATORY COMPLICATIONS|TYPE 1 DIABETES MELLITUS WITH OTH CIRCULATORY COMPLICATIONS
C2832443|T037|S06.4X3S|ICD10CM|EPIDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, SEQUELA|EPIDURAL HEMORRHAGE W LOC OF 1-5 HRS 59 MIN, SEQUELA
C2857565|T037|S72.21XB|ICD10CM|DISPLACED SUBTROCHANTERIC FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPLACED SUBTROCHNT FX R FEMUR, INIT FOR OPN FX TYPE I/2
C4270623|T046|T85.830A|ICD10CM|HEMORRHAGE DUE TO NERVOUS SYSTEM PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|HEMORRHAGE DUE TO NERVOUS SYSTEM PROSTH DEV/GRFT, INIT
C2842086|T191|C50.119|ICD10CM|MALIGNANT NEOPLASM OF CENTRAL PORTION OF UNSPECIFIED FEMALE BREAST|MALIGNANT NEOPLASM OF CENTRAL PORTION OF UNSP FEMALE BREAST
C2882424|T047|I65.29|ICD10CM|OCCLUSION AND STENOSIS OF UNSPECIFIED CAROTID ARTERY|OCCLUSION AND STENOSIS OF UNSPECIFIED CAROTID ARTERY
C3495536|T047|B58.3|DMDICD10|PULMONARY TOXOPLASMOSIS|TOXOPLASMOSE DER LUNGE
C0085315|T047|B58.2|DMDICD10|TOXOPLASMA MENINGOENCEPHALITIS|MENINGOENZEPHALITIS DURCH TOXOPLASMEN
C2832441|T037|S06.4X3A|ICD10CM|EPIDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|EPIDURAL HEMORRHAGE W LOC OF 1-5 HRS 59 MIN, INIT
C2882421|T047|I65.21|ICD10CM|OCCLUSION AND STENOSIS OF RIGHT CAROTID ARTERY|OCCLUSION AND STENOSIS OF RIGHT CAROTID ARTERY
C2882423|T047|I65.23|ICD10CM|OCCLUSION AND STENOSIS OF BILATERAL CAROTID ARTERIES|OCCLUSION AND STENOSIS OF BILATERAL CAROTID ARTERIES
C2882422|T047|I65.22|ICD10CM|OCCLUSION AND STENOSIS OF LEFT CAROTID ARTERY|OCCLUSION AND STENOSIS OF LEFT CAROTID ARTERY
C2874667|T048|F15.929|ICD10CM|OTHER STIMULANT USE, UNSPECIFIED WITH INTOXICATION, UNSPECIFIED|OTHER STIMULANT USE, UNSP WITH INTOXICATION, UNSPECIFIED
C2889239|T047|M05.429|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSP ELBOW
C2874253|T047|E71.528|ICD10CM|OTHER X-LINKED ADRENOLEUKODYSTROPHY|OTHER X-LINKED ADRENOLEUKODYSTROPHY
C0162309|T047|E71.529|ICD10CM|X-LINKED ADRENOLEUKODYSTROPHY, UNSPECIFIED TYPE|X-LINKED ADRENOLEUKODYSTROPHY, UNSPECIFIED TYPE
C4236965|T048|F15.921|ICD10CM|OTHER STIMULANT USE, UNSPECIFIED WITH INTOXICATION DELIRIUM|AMPHETAMINE OR OTHER STIMULANT-INDUCED DELIRIUM
C2874664|T048|F15.920|ICD10CM|OTHER STIMULANT USE, UNSPECIFIED WITH INTOXICATION, UNCOMPLICATED|OTHER STIMULANT USE, UNSP WITH INTOXICATION, UNCOMPLICATED
C2874666|T048|F15.922|ICD10CM|OTHER STIMULANT USE, UNSPECIFIED WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE|OTH STIMULANT USE, UNSP W INTOX W PERCEPTUAL DISTURBANCE
C1527231|T047|E71.522|ICD10CM|ADRENOMYELONEUROPATHY|ADRENOMYELONEUROPATHY
C2889237|T047|M05.421|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT ELBOW|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT ELBOW
C2874249|T047|E71.520|ICD10CM|CHILDHOOD CEREBRAL X-LINKED ADRENOLEUKODYSTROPHY|CHILDHOOD CEREBRAL X-LINKED ADRENOLEUKODYSTROPHY
C2874250|T047|E71.521|ICD10CM|ADOLESCENT X-LINKED ADRENOLEUKODYSTROPHY|ADOLESCENT X-LINKED ADRENOLEUKODYSTROPHY
C2885526|T037|T63.302S|ICD10CM|TOXIC EFFECT OF UNSPECIFIED SPIDER VENOM, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF UNSP SPIDER VENOM, SELF-HARM, SEQUELA
C2865518|T037|S88.011S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT KNEE LEVEL, RIGHT LOWER LEG, SEQUELA|COMPLETE TRAUMATIC AMP AT KNEE LEVEL, R LOW LEG, SEQUELA
C2905787|T037|X81.8XXD|ICD10CM|INTENTIONAL SELF-HARM BY JUMPING OR LYING IN FRONT OF OTHER MOVING OBJECT, SUBSEQUENT ENCOUNTER|SLF-HRM BY JUMPING OR LYING IN FRONT OF MOVING OBJECT, SUBS
C0694505|T047|J99|DMDICD10|RESPIRATORY DISORDERS IN DISEASES CLASSIFIED ELSEWHERE|KRANKHEITEN DER ATEMWEGE BEI ANDERENORTS KLASSIFIZIERTEN KRANKHEITEN
C2976990|T046|I82.4Y1|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF RIGHT PROXIMAL LOWER EXTREMITY|AC EMBLSM AND THOMBOS UNSP DEEP VEINS OF R PROX LOW EXTRM
C2976991|T046|I82.4Y2|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF LEFT PROXIMAL LOWER EXTREMITY|AC EMBLSM AND THOMBOS UNSP DEEP VEINS OF LEFT PROX LOW EXTRM
C2976992|T046|I82.4Y3|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF PROXIMAL LOWER EXTREMITY, BILATERAL|AC EMBLSM AND THOMBOS UNSP DEEP VEINS OF PROX LOW EXTRM, BI
C2859219|T037|S73.033A|ICD10CM|OTHER ANTERIOR SUBLUXATION OF UNSPECIFIED HIP, INITIAL ENCOUNTER|OTHER ANTERIOR SUBLUXATION OF UNSPECIFIED HIP, INIT ENCNTR
C2879415|T037|T46.1X2S|ICD10CM|POISONING BY CALCIUM-CHANNEL BLOCKERS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY CALCIUM-CHANNEL BLOCKERS, SELF-HARM, SEQUELA
C2976993|T046|I82.4Y9|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF UNSPECIFIED PROXIMAL LOWER EXTREMITY|ACUTE EMBLSM AND THOMBOS UNSP DEEP VN UNSP PROX LOW EXTRM
C2833920|T037|S14.121D|ICD10CM|CENTRAL CORD SYNDROME AT C1 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|CENTRAL CORD SYNDROME AT C1, SUBS
C2833919|T037|S14.121A|ICD10CM|CENTRAL CORD SYNDROME AT C1 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|CENTRAL CORD SYNDROME AT C1, INIT
C2874397|T048|F10.259|ICD10CM|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED
C2874395|T048|F10.250|ICD10CM|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|ALCOHOL DEPEND W ALCOH-INDUCE PSYCHOTIC DISORDER W DELUSIONS
C2874396|T048|F10.251|ICD10CM|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|ALCOHOL DEPEND W ALCOH-INDUCE PSYCHOTIC DISORDER W HALLUCIN
C2833921|T037|S14.121S|ICD10CM|CENTRAL CORD SYNDROME AT C1 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|CENTRAL CORD SYNDROME AT C1, SEQUELA
C2901495|T046|M84.653A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, UNSP FEMUR, INIT
C2853966|T191|C84.46|ICD10CM|PERIPHERAL T-CELL LYMPHOMA, NOT CLASSIFIED, INTRAPELVIC LYMPH NODES|PERIPHERAL T-CELL LYMPHOMA, NOT CLASSIFIED, INTRAPELV NODES
C2885884|T037|T63.822A|ICD10CM|TOXIC EFFECT OF CONTACT WITH VENOMOUS TOAD, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CONTACT W VENOMOUS TOAD, SELF-HARM, INIT
C2883811|T037|T50.A12A|ICD10CM|POISONING BY PERTUSSIS VACCINE, INCLUDING COMBINATIONS WITH A PERTUSSIS COMPONENT, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY PERTUSS VACCN, INC COMBIN W PERTUSS, SLF-HRM, INIT
C2853967|T191|C84.47|ICD10CM|PERIPHERAL T-CELL LYMPHOMA, NOT CLASSIFIED, SPLEEN|PERIPHERAL T-CELL LYMPHOMA, NOT CLASSIFIED, SPLEEN
C2853964|T191|C84.44|ICD10CM|PERIPHERAL T-CELL LYMPHOMA, NOT CLASSIFIED, LYMPH NODES OF AXILLA AND UPPER LIMB|PRPH T-CELL LYMPH, NOT CLASS, NODES OF AXILLA AND UPPER LIMB
C2876174|T037|T31.92|ICD10CM|BURNS INVOLVING 90% OR MORE OF BODY SURFACE WITH 20-29% THIRD DEGREE BURNS|BURNS OF 90%/MORE OF BODY SURFC W 20-29% THIRD DEGREE BURNS
C2879413|T037|T46.1X2A|ICD10CM|POISONING BY CALCIUM-CHANNEL BLOCKERS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY CALCIUM-CHANNEL BLOCKERS, SELF-HARM, INIT
C2853965|T191|C84.45|ICD10CM|PERIPHERAL T-CELL LYMPHOMA, NOT CLASSIFIED, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|PRPH T-CELL LYMPH, NOT CLASS, NODES OF ING RGN AND LOW LIMB
C2883813|T037|T50.A12S|ICD10CM|POISONING BY PERTUSSIS VACCINE, INCLUDING COMBINATIONS WITH A PERTUSSIS COMPONENT, INTENTIONAL SELF-HARM, SEQUELA|POISN BY PERTUSS VACCN, INC COMBIN W PERTUSS, SLF-HRM, SQLA
C2853962|T191|C84.42|ICD10CM|PERIPHERAL T-CELL LYMPHOMA, NOT CLASSIFIED, INTRATHORACIC LYMPH NODES|PERIPHERAL T-CELL LYMPHOMA, NOT CLASS, INTRATHORAC NODES
C2877099|T037|T38.4X2S|ICD10CM|POISONING BY ORAL CONTRACEPTIVES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ORAL CONTRACEPTIVES, SELF-HARM, SEQUELA
C2853963|T191|C84.43|ICD10CM|PERIPHERAL T-CELL LYMPHOMA, NOT CLASSIFIED, INTRA-ABDOMINAL LYMPH NODES|PERIPHERAL T-CELL LYMPHOMA, NOT CLASSIFIED, INTRA-ABD NODES
C1456241|T047|G47.429|ICD10CM|NARCOLEPSY IN CONDITIONS CLASSIFIED ELSEWHERE WITHOUT CATAPLEXY|NARCOLEPSY IN CONDITIONS CLASSIFIED ELSEWHERE W/O CATAPLEXY
C4237031|T048|F12.980|ICD10CM|CANNABIS USE, UNSPECIFIED WITH ANXIETY DISORDER|CANNABIS INDUCED ANXIETY DISORDER, WITHOUT USE DISORDER
C1456242|T047|G47.421|ICD10CM|NARCOLEPSY IN CONDITIONS CLASSIFIED ELSEWHERE WITH CATAPLEXY|NARCOLEPSY IN CONDITIONS CLASSIFIED ELSEWHERE WITH CATAPLEXY
C2853961|T191|C84.41|ICD10CM|PERIPHERAL T-CELL LYMPHOMA, NOT CLASSIFIED, LYMPH NODES OF HEAD, FACE, AND NECK|PRPH T-CELL LYMPH, NOT CLASS, NODES OF HEAD, FACE, AND NECK
C2874313|T047|E88.49|ICD10CM|OTHER MITOCHONDRIAL METABOLISM DISORDERS|OTHER MITOCHONDRIAL METABOLISM DISORDERS
C2843277|T037|S48.019A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT UNSPECIFIED SHOULDER JOINT, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION AT UNSP SHOULDER JOINT, INIT
C2845921|T191||ICD10CM|MALIGNANT NEOPLASM OF LEFT ORBIT
C2845920|T191||ICD10CM|MALIGNANT NEOPLASM OF RIGHT ORBIT
C2845919|T191|C69.60|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED ORBIT|MALIGNANT NEOPLASM OF UNSPECIFIED ORBIT
C1456275|T047|E88.40|ICD10CM|MITOCHONDRIAL METABOLISM DISORDER, UNSPECIFIED|MITOCHONDRIAL METABOLISM DISORDER, UNSPECIFIED
C0261612|T067|E884.1|ICD9CM|MELAS SYNDROME|FALL FROM CLIFF
C0261613|T067|E884.2|ICD9CM|MERRF SYNDROME|ACCIDENTAL FALL FROM CHAIR
C2889426|T047|M06.249|ICD10CM|RHEUMATOID BURSITIS, UNSPECIFIED HAND|RHEUMATOID BURSITIS, UNSPECIFIED HAND
C0839988|T047|M86.60|ICD10AM|OTHER CHRONIC OSTEOMYELITIS, UNSPECIFIED SITE|OTHER CHRONIC OSTEOMYELITIS, MULTIPLE SITES
C1397893|T047||ICD10CM|GASTROSTOMY MALFUNCTION
C0695239|T047||ICD10CM|GASTROSTOMY INFECTION
C2888030|T046|K94.21|ICD10CM|GASTROSTOMY HEMORRHAGE|GASTROSTOMY HEMORRHAGE
C0587245|T046|K94.20|ICD10CM|GASTROSTOMY COMPLICATION, UNSPECIFIED|GASTROSTOMY COMPLICATION, UNSPECIFIED
C2889424|T047|M06.241|ICD10CM|RHEUMATOID BURSITIS, RIGHT HAND|RHEUMATOID BURSITIS, RIGHT HAND
C2889425|T047|M06.242|ICD10CM|RHEUMATOID BURSITIS, LEFT HAND|RHEUMATOID BURSITIS, LEFT HAND
C0695241|T046|K94.29|ICD10CM|OTHER COMPLICATIONS OF GASTROSTOMY|OTHER COMPLICATIONS OF GASTROSTOMY
C2874426|T048|F11.129|ICD10CM|OPIOID ABUSE WITH INTOXICATION, UNSPECIFIED|OPIOID ABUSE WITH INTOXICATION, UNSPECIFIED
C2853968|T191|C84.48|ICD10CM|PERIPHERAL T-CELL LYMPHOMA, NOT CLASSIFIED, LYMPH NODES OF MULTIPLE SITES|PERIPHERAL T-CELL LYMPHOMA, NOT CLASSIFIED, NODES MULT SITE
C2858493|T037|S72.424C|ICD10CM|NONDISPLACED FRACTURE OF LATERAL CONDYLE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF LATERAL CONDYLE OF R FEMR, 7THC
C2858492|T037|S72.424B|ICD10CM|NONDISPLACED FRACTURE OF LATERAL CONDYLE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF LATERAL CONDYLE OF R FEMR, 7THB
C0010418|T047|A07.2|DMDICD10|CRYPTOSPORIDIOSIS|KRYPTOSPORIDIOSE
C2874423|T048||ICD10CM|OPIOID ABUSE WITH INTOXICATION, UNCOMPLICATED
C2874425|T048|F11.122|ICD10CM|OPIOID ABUSE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE|OPIOID ABUSE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE
C2885059|T037|T60.3X2A|ICD10CM|TOXIC EFFECT OF HERBICIDES AND FUNGICIDES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF HERBICIDES AND FUNGICIDES, SELF-HARM, INIT
C4267908|T047|E08.3319|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|DIABETES WITH MODERATE NONP RTNOP WITH MACULAR EDEMA, UNSP
C4268002|T047|E09.3591|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|DRUG/CHEM DIAB WITH PROLIF DIAB RTNOP W/O MCLR EDEMA, R EYE
C4268003|T047|E09.3592|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|DRUG/CHEM DIAB WITH PROLIF DIAB RTNOP W/O MCLR EDEMA, L EYE
C4268004|T047|E09.3593|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|DRUG/CHEM DIAB WITH PROLIF DIAB RTNOP WITHOUT MCLR EDEMA, BI
C4267907|T047|E08.3313|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|DIABETES WITH MODERATE NONP RTNOP WITH MACULAR EDEMA, BI
C4267906|T047|E08.3312|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|DIAB WITH MODERATE NONP RTNOP WITH MACULAR EDEMA, LEFT EYE
C4267905|T047|E08.3311|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|DIABETES WITH MODERATE NONP RTNOP WITH MACULAR EDEMA, R EYE
C4268005|T047|E09.3599|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|DRUG/CHEM DIAB WITH PROLIF DIAB RTNOP W/O MCLR EDEMA, UNSP
C2890455|T037|T84.030A|ICD10CM|MECHANICAL LOOSENING OF INTERNAL RIGHT HIP PROSTHETIC JOINT, INITIAL ENCOUNTER|MECH LOOSENING OF INTERNAL RIGHT HIP PROSTHETIC JOINT, INIT
C2901342|T046|M84.575A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, LEFT FOOT, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, LEFT FOOT, INIT
C2837930|T191|C13.1|ICD10CM|MALIGNANT NEOPLASM OF ARYEPIGLOTTIC FOLD, HYPOPHARYNGEAL ASPECT|MALIGNANT NEOPLASM OF INTERARYTENOID FOLD, MARGINAL ZONE
C0496769|T191|C13.0|DMDICD10|MALIGNANT NEOPLASM OF POSTCRICOID REGION|BOESARTIGE NEUBILDUNG: REGIO POSTCRICOIDEA
C0496770|T191|C13.2|DMDICD10|MALIGNANT NEOPLASM OF POSTERIOR WALL OF HYPOPHARYNX|BOESARTIGE NEUBILDUNG: HINTERWAND DES HYPOPHARYNX
C0864862|T191|C13.9|ICD10CM|MALIGNANT NEOPLASM OF HYPOPHARYNX, UNSPECIFIED|MALIGNANT NEOPLASM OF HYPOPHARYNGEAL WALL NOS
C0349039|T191|C13.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF HYPOPHARYNX|BOESARTIGE NEUBILDUNG: HYPOPHARYNX, MEHRERE TEILBEREICHE UEBERLAPPEND
C0300933|T047||ICD10CM|ZYGOMYCOSIS, UNSPECIFIED
C4509281|T047|L97.125|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT THIGH WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OF LEFT THIGH WITH MSL INVL W/O EVD OF NECR
C2888654|T047|L97.124|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT THIGH WITH NECROSIS OF BONE|NON-PRESSURE CHRONIC ULCER OF LEFT THIGH W NECROSIS OF BONE
C0156057|T047|K28.5|DMDICD10|CHRONIC OR UNSPECIFIED GASTROJEJUNAL ULCER WITH PERFORATION|ULCUS PEPTICUM JEJUNI: CHRONISCH ODER NICHT NAEHER BEZEICHNET, MIT PERFORATION
C4509282|T047|L97.126|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT THIGH WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OF LEFT THIGH WITH BONE INVL W/O EVD OF NECR
C2888651|T047|L97.121|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT THIGH LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHRONIC ULCER OF LEFT THIGH LIMITED TO BRKDWN SKIN
C0156048|T047|K28.2|DMDICD10|ACUTE GASTROJEJUNAL ULCER WITH BOTH HEMORRHAGE AND PERFORATION|ULCUS PEPTICUM JEJUNI: AKUT, MIT BLUTUNG UND PERFORATION
C0156045|T047|K28.1|DMDICD10|ACUTE GASTROJEJUNAL ULCER WITH PERFORATION|ULCUS PEPTICUM JEJUNI: AKUT, MIT PERFORATION
C2888652|T047|L97.122|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT THIGH WITH FAT LAYER EXPOSED|NON-PRESSURE CHRONIC ULCER OF LEFT THIGH W FAT LAYER EXPOSED
C2888655|T047|L97.129|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT THIGH WITH UNSPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF LEFT THIGH WITH UNSP SEVERITY
C4509283|T047|L97.128|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT THIGH WITH OTHER SPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF LEFT THIGH WITH OTH SEVERITY
C2861671|T191|D03.30|ICD10CM|MELANOMA IN SITU OF UNSPECIFIED PART OF FACE|MELANOMA IN SITU OF UNSPECIFIED PART OF FACE
C4269431|T037|S02.601S|ICD10CM|FRACTURE OF UNSPECIFIED PART OF BODY OF RIGHT MANDIBLE, SEQUELA|FX UNSPECIFIED PART OF BODY OF RIGHT MANDIBLE, SEQUELA
C2888631|T047|L89.95|ICD10CM|PRESSURE ULCER OF UNSPECIFIED SITE, UNSTAGEABLE|PRESSURE ULCER OF UNSPECIFIED SITE, UNSTAGEABLE
C2888630|T047|L89.94|ICD10CM|PRESSURE ULCER OF UNSPECIFIED SITE, STAGE 4|PRESSURE ULCER OF UNSPECIFIED SITE, STAGE 4
C2888627|T047|L89.93|ICD10CM|PRESSURE ULCER OF UNSPECIFIED SITE, STAGE 3|PRESSURE ULCER OF UNSPECIFIED SITE, STAGE 3
C2888624|T047|L89.92|ICD10CM|PRESSURE ULCER OF UNSPECIFIED SITE, STAGE 2|PRESSURE ULCER OF UNSPECIFIED SITE, STAGE 2
C2861672|T191|D03.39|ICD10CM|MELANOMA IN SITU OF OTHER PARTS OF FACE|MELANOMA IN SITU OF OTHER PARTS OF FACE
C2888618|T047|L89.90|ICD10CM|PRESSURE ULCER OF UNSPECIFIED SITE, UNSPECIFIED STAGE|PRESSURE ULCER OF UNSPECIFIED SITE, UNSPECIFIED STAGE
C4269427|T037|S02.601B|ICD10CM|FRACTURE OF UNSPECIFIED PART OF BODY OF RIGHT MANDIBLE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF UNSPECIFIED PART OF BODY OF RIGHT MANDIBLE, 7THB
C4269426|T037|S02.601A|ICD10CM|FRACTURE OF UNSPECIFIED PART OF BODY OF RIGHT MANDIBLE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF UNSPECIFIED PART OF BODY OF RIGHT MANDIBLE, INIT
C0348492|T047|E76.8|DMDICD10|OTHER DISORDERS OF GLUCOSAMINOGLYCAN METABOLISM|SONSTIGE STOERUNGEN DES GLYKOSAMINOGLYKAN-STOFFWECHSELS
C0348503|T047|E76.9|DMDICD10|GLUCOSAMINOGLYCAN METABOLISM DISORDER, UNSPECIFIED|STOERUNG DES GLYKOSAMINOGLYKAN-STOFFWECHSELS, NICHT NAEHER BEZEICHNET
C0026703|T047|E76.3|DMDICD10|MUCOPOLYSACCHARIDOSIS, UNSPECIFIED|MUKOPOLYSACCHARIDOSE, NICHT NAEHER BEZEICHNET
C0026705|T047|E76.1|DMDICD10|MUCOPOLYSACCHARIDOSIS, TYPE II|MUKOPOLYSACCHARIDOSE, TYP II
C2888460|T047|L89.329|ICD10CM|PRESSURE ULCER OF LEFT BUTTOCK, UNSPECIFIED STAGE|PRESSURE ULCER OF LEFT BUTTOCK, UNSPECIFIED STAGE
C2887643|T047|K22.70|ICD10CM|BARRETT'S ESOPHAGUS WITHOUT DYSPLASIA|BARRETT'S ESOPHAGUS WITHOUT DYSPLASIA
C2888457|T047|L89.324|ICD10CM|PRESSURE ULCER OF LEFT BUTTOCK, STAGE 4|PRESSURE ULCER OF LEFT BUTTOCK, STAGE 4
C2888445|T047||ICD10CM|PRESSURE ULCER OF LEFT BUTTOCK, UNSTAGEABLE
C2888448|T047|L89.321|ICD10CM|PRESSURE ULCER OF LEFT BUTTOCK, STAGE 1|PRESSURE ULCER OF LEFT BUTTOCK, STAGE 1
C2888451|T047|L89.322|ICD10CM|PRESSURE ULCER OF LEFT BUTTOCK, STAGE 2|PRESSURE ULCER OF LEFT BUTTOCK, STAGE 2
C2888454|T047|L89.323|ICD10CM|PRESSURE ULCER OF LEFT BUTTOCK, STAGE 3|PRESSURE ULCER OF LEFT BUTTOCK, STAGE 3
C2838684|T037|S34.125S|ICD10CM|INCOMPLETE LESION OF L5 LEVEL OF LUMBAR SPINAL CORD, SEQUELA|INCOMPLETE LESION OF L5 LEVEL OF LUMBAR SPINAL CORD, SEQUELA
C2901227|T046|M84.542A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, LEFT HAND, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, LEFT HAND, INIT
C4268176|T047|E13.3599|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|OTH DIAB WITH PROLIF DIAB RTNOP WITHOUT MACULAR EDEMA, UNSP
C2875066|T047|G32.0|ICD10CM|SUBACUTE COMBINED DEGENERATION OF SPINAL CORD IN DISEASES CLASSIFIED ELSEWHERE|SCLEROSIS OF SPINAL CORD (COMBINED) (DORSOLATERAL) (POSTEROLATERAL)
C2865539|T037|S88.029S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT KNEE LEVEL, UNSPECIFIED LOWER LEG, SEQUELA|PARTIAL TRAUMATIC AMP AT KNEE LEVEL, UNSP LOWER LEG, SEQUELA
C4268173|T047|E13.3591|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|OTH DIAB WITH PROLIF DIAB RTNOP WITHOUT MACULAR EDEMA, R EYE
C4268175|T047|E13.3593|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|OTH DIAB WITH PROLIF DIAB RTNOP WITHOUT MACULAR EDEMA, BI
C4268174|T047|E13.3592|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|OTH DIAB WITH PROLIF DIAB RTNOP WITHOUT MACULAR EDEMA, L EYE
C2891282|T037|T86.49|ICD10CM|OTHER COMPLICATIONS OF LIVER TRANSPLANT|OTHER COMPLICATIONS OF LIVER TRANSPLANT
C2858012|T037|S72.346C|ICD10CM|NONDISPLACED SPIRAL FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP SPIRAL FX SHAFT OF UNSP FEMR, 7THC
C2833584|T037|S12.600A|ICD10CM|UNSPECIFIED DISPLACED FRACTURE OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP DISP FX OF SEVENTH CERVICAL VERTEBRA, INIT FOR CLOS FX
C1444565|T046|R09.2|ICD10CM|RESPIRATORY ARREST|CARDIORESPIRATORY FAILURE
C2865537|T037|S88.029A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT KNEE LEVEL, UNSPECIFIED LOWER LEG, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP AT KNEE LEVEL, UNSP LOWER LEG, INIT
C0400969|T046|T86.42|ICD10CM|LIVER TRANSPLANT FAILURE|LIVER TRANSPLANT FAILURE
C0400968|T046|T86.41|ICD10CM|LIVER TRANSPLANT REJECTION|LIVER TRANSPLANT REJECTION
C2833779|T037|S14.102A|ICD10CM|UNSPECIFIED INJURY AT C2 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY AT C2 LEVEL OF CERVICAL SPINAL CORD, INIT ENCNTR
C2865538|T037|S88.029D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT KNEE LEVEL, UNSPECIFIED LOWER LEG, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMP AT KNEE LEVEL, UNSP LOWER LEG, SUBS
C2833851|T037|S14.102D|ICD10CM|UNSPECIFIED INJURY AT C2 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY AT C2 LEVEL OF CERVICAL SPINAL CORD, SUBS ENCNTR
C2882503|T047|I69.149|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING UNSPECIFIED SIDE|MONOPLG LOW LMB FOLLOWING NTRM INTCRBL HEMOR AFF UNSP SIDE
C2889491|T047|M06.879|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, UNSPECIFIED ANKLE AND FOOT|OTH RHEUMATOID ARTHRITIS, UNSPECIFIED ANKLE AND FOOT
C2882499|T047|I69.141|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING RIGHT DOMINANT SIDE|MONOPLG LOW LMB FOL NTRM INTCRBL HEMOR AFF RIGHT DOM SIDE
C2882501|T047|I69.143|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING RIGHT NON-DOMINANT SIDE|MONOPLG LOW LMB FOL NTRM INTCRBL HEMOR AFF RIGHT NONDOM SIDE
C2882500|T047|I69.142|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING LEFT DOMINANT SIDE|MONOPLG LOW LMB FOL NTRM INTCRBL HEMOR AFF LEFT DOM SIDE
C2882502|T047|I69.144|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING LEFT NON-DOMINANT SIDE|MONOPLG LOW LMB FOL NTRM INTCRBL HEMOR AFF LEFT NONDOM SIDE
C2873867|T047|E05.10|ICD10CM|THYROTOXICOSIS WITH TOXIC SINGLE THYROID NODULE WITHOUT THYROTOXIC CRISIS OR STORM|THYROTXCOSIS W TOXIC SING THYROID NODULE W/O THYROTXC CRISIS
C0154141|T047|E05.11|ICD10CM|THYROTOXICOSIS WITH TOXIC SINGLE THYROID NODULE WITH THYROTOXIC CRISIS OR STORM|THYROTOXICOSIS WITH TOXIC SINGLE THYROID NODULE WITH THYROTOXIC CRISIS OR STORM
C0840039|T046|M87.39|ICD10CM|OTHER SECONDARY OSTEONECROSIS, MULTIPLE SITES|OTHER SECONDARY OSTEONECROSIS, MULTIPLE SITES
C2875116|T047|G40.419|ICD10CM|OTHER GENERALIZED EPILEPSY AND EPILEPTIC SYNDROMES, INTRACTABLE, WITHOUT STATUS EPILEPTICUS|OTH GENERALIZED EPILEPSY, INTRACTABLE, W/O STAT EPI
C2858903|T037|S72.464B|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP SUPRCNDL FX W INTRCNDL EXTN LOW END R FEMR, 7THB
C1387047|T048||ICD10CM|BORDERLINE PERSONALITY DISORDER
C2886880|T037|T81.502S|ICD10CM|UNSPECIFIED COMPLICATION OF FOREIGN BODY ACCIDENTALLY LEFT IN BODY FOLLOWING KIDNEY DIALYSIS, SEQUELA|UNSP COMP OF FB ACC LEFT IN BODY FOL KIDNEY DIALYSIS, SQLA
C1704373|T048||ICD10CM|OBSESSIVE-COMPULSIVE PERSONALITY DISORDER
C2832309|T037|S06.361A|ICD10CM|TRAUMATIC HEMORRHAGE OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|TRAUM HEMOR CEREB, W LOC OF 30 MINUTES OR LESS, INIT
C2843344|T037|S48.929S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED SHOULDER AND UPPER ARM, LEVEL UNSPECIFIED, SEQUELA|PARTIAL TRAUM AMP OF UNSP SHLDR/UP ARM, LEVEL UNSP, SEQUELA
C2896477|T046|M80.00XA|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, UNSPECIFIED SITE, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, UNSP SITE, INIT
C2901896|T047|M86.529|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED HUMERUS|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, UNSP HUMERUS
C2886878|T037|T81.502A|ICD10CM|UNSPECIFIED COMPLICATION OF FOREIGN BODY ACCIDENTALLY LEFT IN BODY FOLLOWING KIDNEY DIALYSIS, INITIAL ENCOUNTER|UNSP COMP OF FB ACC LEFT IN BODY FOL KIDNEY DIALYSIS, INIT
C2832311|T037|S06.361S|ICD10CM|TRAUMATIC HEMORRHAGE OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|TRAUM HEMOR CEREB, W LOC OF 30 MINUTES OR LESS, SEQUELA
C2901894|T047|M86.521|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, RIGHT HUMERUS|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, RIGHT HUMERUS
C2895319|T037|M48.52XA|ICD10CM|COLLAPSED VERTEBRA, NOT ELSEWHERE CLASSIFIED, CERVICAL REGION, INITIAL ENCOUNTER FOR FRACTURE|COLLAPSED VERTEBRA, NEC, CERVICAL REGION, INIT
C2887465|T047|J45.909|ICD10CM|UNSPECIFIED ASTHMA, UNCOMPLICATED|UNSPECIFIED ASTHMA, UNCOMPLICATED
C2835319|T037|S22.048A|ICD10CM|OTHER FRACTURE OF FOURTH THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF FOURTH THORACIC VERTEBRA, INIT FOR CLOS FX
C2835320|T037|S22.048B|ICD10CM|OTHER FRACTURE OF FOURTH THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF FOURTH THORACIC VERTEBRA, INIT FOR OPN FX
C2887464|T047|J45.902|ICD10CM|UNSPECIFIED ASTHMA WITH STATUS ASTHMATICUS|UNSPECIFIED ASTHMA WITH STATUS ASTHMATICUS
C2887463|T047|J45.901|ICD10CM|UNSPECIFIED ASTHMA WITH (ACUTE) EXACERBATION|UNSPECIFIED ASTHMA WITH (ACUTE) EXACERBATION
C2835762|T037|S24.102S|ICD10CM|UNSPECIFIED INJURY AT T2-T6 LEVEL OF THORACIC SPINAL CORD, SEQUELA|UNSP INJURY AT T2-T6 LEVEL OF THORACIC SPINAL CORD, SEQUELA
C2874081|T047|E11.311|ICD10CM|TYPE 2 DIABETES MELLITUS WITH UNSPECIFIED DIABETIC RETINOPATHY WITH MACULAR EDEMA|TYPE 2 DIABETES W UNSP DIABETIC RETINOPATHY W MACULAR EDEMA
C2874082|T047|E11.319|ICD10CM|TYPE 2 DIABETES MELLITUS WITH UNSPECIFIED DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA|TYPE 2 DIABETES W UNSP DIABETIC RTNOP W/O MACULAR EDEMA
C2901423|T046|M84.632A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, LEFT ULNA, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, LEFT ULNA, INIT FOR FX
C2882345|T047|I63.12|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF BASILAR ARTERY|CEREBRAL INFARCTION DUE TO EMBOLISM OF BASILAR ARTERY
C2882340|T047|I63.10|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF UNSPECIFIED PRECEREBRAL ARTERY|CEREBRAL INFARCTION DUE TO EMBOLISM OF UNSP PRECERB ARTERY
C2882852|T047|I70.491|ICD10CM|OTHER ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES, RIGHT LEG|OTH ATHSCL AUTOLOGOUS VEIN BYPASS OF THE EXTRM, RIGHT LEG
C2902449|T047|M90.571|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, RIGHT ANKLE AND FOOT|OSTEONECROSIS IN DISEASES CLASSD ELSWHR, RIGHT ANK/FT
C2882854|T047|I70.493|ICD10CM|OTHER ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES, BILATERAL LEGS|OTH ATHSCL AUTOL VEIN BYPASS OF THE EXTRM, BILATERAL LEGS
C2882853|T047|I70.492|ICD10CM|OTHER ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES, LEFT LEG|OTH ATHSCL AUTOLOGOUS VEIN BYPASS OF THE EXTRM, LEFT LEG
C0473224|T047|M83.4|DMDICD10|ALUMINUM BONE DISEASE|ALUMINIUMOSTEOPATHIE
C2882350|T047|I63.19|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF OTHER PRECEREBRAL ARTERY|CEREBRAL INFARCTION DUE TO EMBOLISM OF PRECEREBRAL ARTERY
C2882856|T047|I70.499|ICD10CM|OTHER ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES, UNSPECIFIED EXTREMITY|OTH ATHSCL AUTOL VEIN BYPASS OF THE EXTRM, UNSP EXTREMITY
C2882855|T047|I70.498|ICD10CM|OTHER ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES, OTHER EXTREMITY|OTH ATHSCL AUTOL VEIN BYPASS OF THE EXTRM, OTH EXTREMITY
C0410446|T047|M83.0|DMDICD10|PUERPERAL OSTEOMALACIA|OSTEOMALAZIE IM WOCHENBETT
C0451874|T047|M83.1|DMDICD10|SENILE OSTEOMALACIA|SENILE OSTEOMALAZIE
C2876893|T037|T37.4X2A|ICD10CM|POISONING BY ANTHELMINTHICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ANTHELMINTHICS, INTENTIONAL SELF-HARM, INIT
C4290162|T047|I70.45|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF OTHER EXTREMITY WITH ULCERATION|ANY CONDITION CLASSIFIABLE TO I70.418, I70.428, AND I70.438
C2876920|T037|T37.5X2S|ICD10CM|POISONING BY ANTIVIRAL DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ANTIVIRAL DRUGS, INTENTIONAL SELF-HARM, SEQUELA
C2838480|T037|S32.692B|ICD10CM|OTHER SPECIFIED FRACTURE OF LEFT ISCHIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF LEFT ISCHIUM, INIT ENCNTR FOR OPEN FRACTURE
C0477970|T019|Q03.8|DMDICD10|OTHER CONGENITAL HYDROCEPHALUS|SONSTIGER ANGEBORENER HYDROZEPHALUS
C0020256|T019|Q03|DMDICD10|CONGENITAL HYDROCEPHALUS, UNSPECIFIED|ANGEBORENER HYDROZEPHALUS
C0266476|T019||ICD10CM|MALFORMATIONS OF AQUEDUCT OF SYLVIUS
C0010964|T047|Q03.1|DMDICD10|ATRESIA OF FORAMINA OF MAGENDIE AND LUSCHKA|ATRESIE DER APERTURA MEDIANA [FORAMEN MAGENDII] ODER DER APERTURAE LATERALES [FORAMINA LUSCHKAE] DES VIERTEN VENTRIKELS
C2876918|T037|T37.5X2A|ICD10CM|POISONING BY ANTIVIRAL DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ANTIVIRAL DRUGS, INTENTIONAL SELF-HARM, INIT
C2833293|T037|S12.151A|ICD10CM|OTHER TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH TRAUM NONDISP SPONDYLOLYSIS OF SECOND CERVCAL VERT, INIT
C2833294|T037|S12.151B|ICD10CM|OTHER TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH TRAUM NONDISP SPONDYLOLYSIS OF 2ND CERVCAL VERT, 7THB
C2887833|T047||ICD10CM|OTHER ULCERATIVE COLITIS WITH INTESTINAL OBSTRUCTION
C2887834|T047||ICD10CM|OTHER ULCERATIVE COLITIS WITH FISTULA
C2873806|T046|D69.3|ICD10CM|IMMUNE THROMBOCYTOPENIC PURPURA|HEMORRHAGIC (THROMBOCYTOPENIC) PURPURA
C2887832|T047||ICD10CM|OTHER ULCERATIVE COLITIS WITH RECTAL BLEEDING
C2887835|T047||ICD10CM|OTHER ULCERATIVE COLITIS WITH ABSCESS
C0040034|T047|D69.6|DMDICD10|THROMBOCYTOPENIA, UNSPECIFIED|THROMBOZYTOPENIE, NICHT NAEHER BEZEICHNET
C0019087|T047|D69.9|DMDICD10|HEMORRHAGIC CONDITION, UNSPECIFIED|HAEMORRHAGISCHE DIATHESE, NICHT NAEHER BEZEICHNET
C0340804|T047||ICD10CM|OTHER SPECIFIED HEMORRHAGIC CONDITIONS
C2887836|T047|K51.818|ICD10CM|OTHER ULCERATIVE COLITIS WITH OTHER COMPLICATION|OTHER ULCERATIVE COLITIS WITH OTHER COMPLICATION
C2887837|T047|K51.819|ICD10CM|OTHER ULCERATIVE COLITIS WITH UNSPECIFIED COMPLICATIONS|OTHER ULCERATIVE COLITIS WITH UNSPECIFIED COMPLICATIONS
C2832533|T037|S06.6X6A|ICD10CM|TRAUMATIC SUBARACHNOID HEMORRHAGE WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|TRAUM SUBRAC HEM W LOC >24 HR W/O RET CONSC W SURV, INIT
C2831560|T037|S02.66XB|ICD10CM|FRACTURE OF SYMPHYSIS OF MANDIBLE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF SYMPHYSIS OF MANDIBLE, INIT FOR OPN FX
C2831559|T037|S02.66XA|ICD10CM|FRACTURE OF SYMPHYSIS OF MANDIBLE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF SYMPHYSIS OF MANDIBLE, INIT FOR CLOS FX
C2832535|T037|S06.6X6S|ICD10CM|TRAUMATIC SUBARACHNOID HEMORRHAGE WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|TRAUM SUBRAC HEM W LOC >24 HR W/O RET CONSC W SURV, SEQUELA
C2831564|T037|S02.66XS|ICD10CM|FRACTURE OF SYMPHYSIS OF MANDIBLE, SEQUELA|FRACTURE OF SYMPHYSIS OF MANDIBLE, SEQUELA
C4270205|T046|T83.022A|ICD10CM|DISPLACEMENT OF NEPHROSTOMY CATHETER, INITIAL ENCOUNTER|DISPLACEMENT OF NEPHROSTOMY CATHETER, INITIAL ENCOUNTER
C2874530|T048|F13.220|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH INTOXICATION, UNCOMPLICATED|SEDATV/HYP/ANXIOLYTC DEPENDENCE W INTOXICATION, UNCOMP
C2874531|T048|F13.221|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH INTOXICATION DELIRIUM|SEDATV/HYP/ANXIOLYTC DEPENDENCE W INTOXICATION DELIRIUM
C0494788|T047|K73.1|DMDICD10|CHRONIC LOBULAR HEPATITIS, NOT ELSEWHERE CLASSIFIED|CHRONISCHE LOBULAERE HEPATITIS, ANDERENORTS NICHT KLASSIFIZIERT
C0494787|T047|K73.0|DMDICD10|CHRONIC PERSISTENT HEPATITIS, NOT ELSEWHERE CLASSIFIED|CHRONISCHE PERSISTIERENDE HEPATITIS, ANDERENORTS NICHT KLASSIFIZIERT
C2874532|T048|F13.22|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH INTOXICATION, UNSPECIFIED|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH INTOXICATION
C0019189|T047|K73.9|DMDICD10|CHRONIC HEPATITIS, UNSPECIFIED|CHRONISCHE HEPATITIS, NICHT NAEHER BEZEICHNET
C0494790|T047|K73.8|DMDICD10|OTHER CHRONIC HEPATITIS, NOT ELSEWHERE CLASSIFIED|SONSTIGE CHRONISCHE HEPATITIS, ANDERENORTS NICHT KLASSIFIZIERT
C2858251|T037|S72.392A|ICD10CM|OTHER FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF SHAFT OF LEFT FEMUR, INIT FOR CLOS FX
C2858253|T037|S72.392C|ICD10CM|OTHER FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|OTH FX SHAFT OF LEFT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2858252|T037|S72.392B|ICD10CM|OTHER FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|OTH FX SHAFT OF LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C0025162|T047||ICD10CM|TOXIC MEGACOLON
C4267961|T047|E09.3299|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|DRUG/CHEM DIAB WITH MILD NONP RTNOP WITHOUT MCLR EDEMA, UNSP
C2890871|T037|T84.623A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL FIXATION DEVICE OF LEFT TIBIA, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INT FIX OF LEFT TIBIA, INIT
C2833443|T037|S12.391B|ICD10CM|OTHER NONDISPLACED FRACTURE OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH NONDISP FX OF FOURTH CERVICAL VERTEBRA, INIT FOR OPN FX
C2879846|T037|T47.7X2A|ICD10CM|POISONING BY EMETICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY EMETICS, INTENTIONAL SELF-HARM, INIT ENCNTR
C2833442|T037|S12.391A|ICD10CM|OTHER NONDISPLACED FRACTURE OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH NONDISP FX OF FOURTH CERVICAL VERTEBRA, INIT FOR CLOS FX
C4267960|T047|E09.3293|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|DRUG/CHEM DIAB WITH MILD NONP RTNOP WITHOUT MCLR EDEMA, BI
C4267959|T047|E09.3292|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|DRUG/CHEM DIAB WITH MILD NONP RTNOP W/O MCLR EDEMA, L EYE
C4267958|T047|E09.3291|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|DRUG/CHEM DIAB WITH MILD NONP RTNOP W/O MCLR EDEMA, R EYE
C4290132|T047|I10|ICD10CM|ESSENTIAL (PRIMARY) HYPERTENSION|HYPERTENSION (ARTERIAL) (BENIGN) (ESSENTIAL) (MALIGNANT) (PRIMARY) (SYSTEMIC)
C0837507|T047|M05.00|ICD10AM|FELTY'S SYNDROME, UNSPECIFIED SITE|FELTY'S SYNDROME, MULTIPLE SITES
C2845887|T191|C63.8|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF MALE GENITAL ORGANS|PRIMARY MALIGNANT NEOPLASM OF TWO OR MORE CONTIGUOUS SITES OF MALE GENITAL ORGANS WHOSE POINT OF ORIGIN CANNOT BE DETERMINED
C2845888|T191|C63.9|ICD10CM|MALIGNANT NEOPLASM OF MALE GENITAL ORGAN, UNSPECIFIED|MALIGNANT NEOPLASM OF MALE GENITOURINARY TRACT NOS
C0348368|T191|C63.7|DMDICD10|MALIGNANT NEOPLASM OF OTHER SPECIFIED MALE GENITAL ORGANS|BOESARTIGE NEUBILDUNG: SONSTIGE NAEHER BEZEICHNETE MAENNLICHE GENITALORGANE
C0864963|T191|C63.2|ICD10CM|MALIGNANT NEOPLASM OF SCROTUM|MALIGNANT NEOPLASM OF SKIN OF SCROTUM
C2901976|T046|M87.071|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF RIGHT ANKLE|IDIOPATHIC ASEPTIC NECROSIS OF RIGHT ANKLE
C2901978|T046|M87.073|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED ANKLE|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED ANKLE
C2901977|T046|M87.072|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF LEFT ANKLE|IDIOPATHIC ASEPTIC NECROSIS OF LEFT ANKLE
C2901980|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF LEFT FOOT
C2901979|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF RIGHT FOOT
C2901982|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF RIGHT TOE(S)
C2901981|T046|M87.076|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED FOOT|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED FOOT
C2901984|T046|M87.079|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED TOE(S)|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED TOE(S)
C2901983|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF LEFT TOE(S)
C2865581|T037|S88.921A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT LOWER LEG, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF R LOW LEG, LEVEL UNSP, INIT
C2865582|T037|S88.921D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT LOWER LEG, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF R LOW LEG, LEVEL UNSP, SUBS
C2889167|T047|M05.212|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT SHOULDER|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF L SHOULDER
C2889166|T047|M05.211|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT SHOULDER|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF R SHOULDER
C2889340|T047|M05.741|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT HAND WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRITIS W RHEU FACTOR OF R HAND W/O ORG/SYS INVOLV
C2889341|T047|M05.742|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HAND WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRITIS W RHEU FACTOR OF LEFT HAND W/O ORG/SYS INVOLV
C2865583|T037|S88.921S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT LOWER LEG, LEVEL UNSPECIFIED, SEQUELA|PARTIAL TRAUMATIC AMP OF R LOW LEG, LEVEL UNSP, SEQUELA
C2889168|T047|M05.219|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER
C2883533|T037|T50.0X2A|ICD10CM|POISONING BY MINERALOCORTICOIDS AND THEIR ANTAGONISTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY MINERALOCORTICOIDS AND ANTAG, SELF-HARM, INIT
C2889342|T047|M05.749|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED HAND WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRITIS W RHEU FACTOR OF UNSP HAND W/O ORG/SYS INVOLV
C2838465|T037|S32.616B|ICD10CM|NONDISPLACED AVULSION FRACTURE OF UNSPECIFIED ISCHIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP AVULSION FRACTURE OF UNSP ISCHIUM, INIT FOR OPN FX
C2838464|T037|S32.616A|ICD10CM|NONDISPLACED AVULSION FRACTURE OF UNSPECIFIED ISCHIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED AVULSION FRACTURE OF UNSP ISCHIUM, INIT
C2837603|T037|S32.042A|ICD10CM|UNSTABLE BURST FRACTURE OF FOURTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSTABLE BURST FRACTURE OF FOURTH LUMBAR VERTEBRA, INIT
C2833599|T037|S12.630A|ICD10CM|UNSPECIFIED TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP TRAUM DISPL SPONDYLOLYSIS OF SEVENTH CERVCAL VERT, INIT
C2833600|T037|S12.630B|ICD10CM|UNSPECIFIED TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP TRAUM DISPL SPONDYLOLYSIS OF 7TH CERVCAL VERT, 7THB
C2874629|T048|F15.121|ICD10CM|OTHER STIMULANT ABUSE WITH INTOXICATION DELIRIUM|OTHER STIMULANT ABUSE WITH INTOXICATION DELIRIUM
C2874628|T048|F15.120|ICD10CM|OTHER STIMULANT ABUSE WITH INTOXICATION, UNCOMPLICATED|OTHER STIMULANT ABUSE WITH INTOXICATION, UNCOMPLICATED
C4268243|T048|F15.122|ICD10CM|OTHER STIMULANT ABUSE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE|AMPHETAMINE OR OTHER STIMULANT USE DISORDER, MILD, WITH AMPHETAMINE OR OTHER STIMULANT INTOXICATION, WITH PERCEPTUAL DISTURBANCES
C2887303|T047|I87.319|ICD10CM|CHRONIC VENOUS HYPERTENSION (IDIOPATHIC) WITH ULCER OF UNSPECIFIED LOWER EXTREMITY|CHRONIC VENOUS HYPERTENSION W ULCER OF UNSP LOW EXTRM
C4268244|T048|F15.129|ICD10CM|OTHER STIMULANT ABUSE WITH INTOXICATION, UNSPECIFIED|AMPHETAMINE OR OTHER STIMULANT USE DISORDER, MILD, WITH AMPHETAMINE OR OTHER STIMULANT INTOXICATION, WITHOUT PERCEPTUAL DISTURBANCES
C2882386|T047|I63.421|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF RIGHT ANTERIOR CEREBRAL ARTERY|CEREBRAL INFRC DUE TO EMBOLISM OF RIGHT ANT CEREBRAL ARTERY
C2882387|T047|I63.422|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF LEFT ANTERIOR CEREBRAL ARTERY|CEREBRAL INFRC DUE TO EMBOLISM OF LEFT ANT CEREBRAL ARTERY
C4268486|T047|I63.423|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF BILATERAL ANTERIOR CEREBRAL ARTERIES|CEREBRAL INFRC DUE TO EMBOLISM OF BI ANT CEREBRAL ARTERIES
C2869839|T037|S98.212D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF TWO OR MORE LEFT LESSER TOES, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMP OF TWO OR MORE LEFT LESSER TOES, SUBS
C2869840|T037|S98.212S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF TWO OR MORE LEFT LESSER TOES, SEQUELA|COMPLETE TRAUM AMP OF TWO OR MORE LEFT LESSER TOES, SEQUELA
C2856065|T037|S68.625S|ICD10CM|PARTIAL TRAUMATIC TRANSPHALANGEAL AMPUTATION OF LEFT RING FINGER, SEQUELA|PARTIAL TRAUMATIC TRNSPHAL AMPUTATION OF L RNG FNGR, SEQUELA
C2883113|T046|I82.491|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF OTHER SPECIFIED DEEP VEIN OF RIGHT LOWER EXTREMITY|ACUTE EMBOLISM AND THROMBOSIS OF DEEP VEIN OF R LOW EXTREM
C0153384|T191|C09.0|DMDICD10|MALIGNANT NEOPLASM OF TONSILLAR FOSSA|BOESARTIGE NEUBILDUNG: FOSSA TONSILLARIS
C0153385|T191|C09.1|DMDICD10|MALIGNANT NEOPLASM OF TONSILLAR PILLAR (ANTERIOR) (POSTERIOR)|BOESARTIGE NEUBILDUNG: GAUMENBOGEN (VORDERER) (HINTERER)
C2873810|T046|D70.1|ICD10CM|AGRANULOCYTOSIS SECONDARY TO CANCER CHEMOTHERAPY|AGRANULOCYTOSIS SECONDARY TO CANCER CHEMOTHERAPY
C2845931|T191|C72.22|ICD10CM|MALIGNANT NEOPLASM OF LEFT OLFACTORY NERVE|MALIGNANT NEOPLASM OF LEFT OLFACTORY NERVE
C2845930|T191|C72.21|ICD10CM|MALIGNANT NEOPLASM OF RIGHT OLFACTORY NERVE|MALIGNANT NEOPLASM OF RIGHT OLFACTORY NERVE
C3263992|T047|G40.A09|ICD10CM|ABSENCE EPILEPTIC SYNDROME, NOT INTRACTABLE, WITHOUT STATUS EPILEPTICUS|ABSENCE EPILEPTIC SYNDROME, NOT INTRACTABLE, W/O STAT EPI
C2834054|T037|S14.156S|ICD10CM|OTHER INCOMPLETE LESION AT C6 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|OTH INCOMPLETE LESION AT C6, SEQUELA
C2834053|T037|S14.156D|ICD10CM|OTHER INCOMPLETE LESION AT C6 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|OTH INCOMPLETE LESION AT C6, SUBS
C2858920|T037|S72.465B|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP SUPRCNDL FX W INTRCNDL EXTN LOW END L FEMR, 7THB
C2835799|T037|S24.131S|ICD10CM|ANTERIOR CORD SYNDROME AT T1 LEVEL OF THORACIC SPINAL CORD, SEQUELA|ANTERIOR CORD SYNDROME AT T1, SEQUELA
C2834052|T037|S14.156A|ICD10CM|OTHER INCOMPLETE LESION AT C6 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|OTH INCOMPLETE LESION AT C6, INIT
C2858919|T037|S72.465A|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP SUPRCNDL FX W INTRCNDL EXTN LOWER END L FEMUR, INIT
C2842100|T191|C50.319|ICD10CM|MALIGNANT NEOPLASM OF LOWER-INNER QUADRANT OF UNSPECIFIED FEMALE BREAST|MALIG NEOPLASM OF LOWER-INNER QUADRANT OF UNSP FEMALE BREAST
C4269368|T037|S02.401S|ICD10CM|MAXILLARY FRACTURE, UNSPECIFIED SIDE, SEQUELA|MAXILLARY FRACTURE, UNSPECIFIED SIDE, SEQUELA
C4268802|T046|M84.758A|ICD10CM|COMPLETE OBLIQUE ATYPICAL FEMORAL FRACTURE, LEFT LEG, INITIAL ENCOUNTER FOR FRACTURE|COMPLETE OBLIQUE ATYPICAL FEMORAL FRACTURE, LEFT LEG, INIT
C2875106|T047|G40.309|ICD10CM|GENERALIZED IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES, NOT INTRACTABLE, WITHOUT STATUS EPILEPTICUS|GEN IDIOPATHIC EPILEPSY, NOT INTRACTABLE, W/O STAT EPI
C2873812|T047|D70.8|ICD10CM|OTHER NEUTROPENIA|OTHER NEUTROPENIA
C2875105|T047|G40.301|ICD10CM|GENERALIZED IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES, NOT INTRACTABLE, WITH STATUS EPILEPTICUS|GENERALIZED IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES, NOT INTRACTABLE, WITH STATUS EPILEPTICUS
C2885373|T037|T63.042A|ICD10CM|TOXIC EFFECT OF COBRA VENOM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF COBRA VENOM, INTENTIONAL SELF-HARM, INIT
C2856092|T037|S68.712S|ICD10CM|COMPLETE TRAUMATIC TRANSMETACARPAL AMPUTATION OF LEFT HAND, SEQUELA|COMPLETE TRAUMATIC TRANSMETCRPL AMP OF LEFT HAND, SEQUELA
C2887759|T047|K50.019|ICD10CM|CROHN'S DISEASE OF SMALL INTESTINE WITH UNSPECIFIED COMPLICATIONS|CROHN'S DISEASE OF SMALL INTESTINE WITH UNSP COMPLICATIONS
C0271923|T047|D60.0|DMDICD10|CHRONIC ACQUIRED PURE RED CELL APLASIA|CHRONISCHE ERWORBENE ISOLIERTE APLASTISCHE ANAEMIE
C2887758|T047|K50.018|ICD10CM|CROHN'S DISEASE OF SMALL INTESTINE WITH OTHER COMPLICATION|CROHN'S DISEASE OF SMALL INTESTINE WITH OTHER COMPLICATION
C0496902|T191|D35.3|DMDICD10|BENIGN NEOPLASM OF CRANIOPHARYNGEAL DUCT|GUTARTIGE NEUBILDUNG: DUCTUS CRANIOPHARYNGEALIS
C2856090|T037|S68.712A|ICD10CM|COMPLETE TRAUMATIC TRANSMETACARPAL AMPUTATION OF LEFT HAND, INITIAL ENCOUNTER|COMPLETE TRAUMATIC TRANSMETCRPL AMP OF LEFT HAND, INIT
C0261227|T067|E830.1|ICD9CM|WILSON'S DISEASE|BOAT ACC W SUBMERS-POWER
C0261226|T067|E830.0|ICD9CM|DISORDER OF COPPER METABOLISM, UNSPECIFIED|BOAT ACC W SUBMERS-UNPOW
C2882973|T047|I70.701|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, RIGHT LEG|UNSP ATHSCL TYPE OF BYPASS OF THE EXTREMITIES, RIGHT LEG
C2882975|T047|I70.703|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, BILATERAL LEGS|UNSP ATHSCL TYPE OF BYPASS OF THE EXTRM, BILATERAL LEGS
C2882974|T047|I70.702|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, LEFT LEG|UNSP ATHSCL TYPE OF BYPASS OF THE EXTREMITIES, LEFT LEG
C2874298|T047|E83.09|ICD10CM|OTHER DISORDERS OF COPPER METABOLISM|OTHER DISORDERS OF COPPER METABOLISM
C2882977|T047|I70.709|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, UNSPECIFIED EXTREMITY|UNSP ATHSCL TYPE OF BYPASS OF THE EXTRM, UNSP EXTREMITY
C2882976|T047|I70.708|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, OTHER EXTREMITY|UNSP ATHSCL TYPE OF BYPASS OF THE EXTREMITIES, OTH EXTREMITY
C2860171|T037|S79.122A|ICD10CM|SALTER-HARRIS TYPE II PHYSEAL FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SLTR-HARIS TYPE II PHYSEAL FX LOWER END OF LEFT FEMUR, INIT
C2888505|T047|L89.513|ICD10CM|PRESSURE ULCER OF RIGHT ANKLE, STAGE 3|PRESSURE ULCER OF RIGHT ANKLE, STAGE 3
C2888502|T047|L89.512|ICD10CM|PRESSURE ULCER OF RIGHT ANKLE, STAGE 2|PRESSURE ULCER OF RIGHT ANKLE, STAGE 2
C2888499|T047|L89.511|ICD10CM|PRESSURE ULCER OF RIGHT ANKLE, STAGE 1|PRESSURE ULCER OF RIGHT ANKLE, STAGE 1
C2888496|T047||ICD10CM|PRESSURE ULCER OF RIGHT ANKLE, UNSTAGEABLE
C2888508|T047|L89.514|ICD10CM|PRESSURE ULCER OF RIGHT ANKLE, STAGE 4|PRESSURE ULCER OF RIGHT ANKLE, STAGE 4
C0153916|T191|C94.81|ICD10CM|OTHER SPECIFIED LEUKEMIAS, IN REMISSION|OTHER SPECIFIED LEUKEMIAS, IN REMISSION
C2861643|T191|C94.80|ICD10CM|OTHER SPECIFIED LEUKEMIAS NOT HAVING ACHIEVED REMISSION|OTHER SPECIFIED LEUKEMIAS NOT HAVING ACHIEVED REMISSION
C2888511|T047|L89.519|ICD10CM|PRESSURE ULCER OF RIGHT ANKLE, UNSPECIFIED STAGE|PRESSURE ULCER OF RIGHT ANKLE, UNSPECIFIED STAGE
C2349303|T191|C94.82|ICD10CM|OTHER SPECIFIED LEUKEMIAS, IN RELAPSE|OTHER SPECIFIED LEUKEMIAS, IN RELAPSE
C0348946|T047|E74.4|DMDICD10|DISORDERS OF PYRUVATE METABOLISM AND GLUCONEOGENESIS|STOERUNGEN DES PYRUVATSTOFFWECHSELS UND DER GLUKONEOGENESE
C2837737|T037|S32.131B|ICD10CM|MINIMALLY DISPLACED ZONE III FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|MINIMALLY DISPLACED ZONE III FX SACRUM, INIT FOR OPN FX
C2901918|T047|M86.629|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, UNSPECIFIED  HUMERUS|OTHER CHRONIC OSTEOMYELITIS, UNSPECIFIED HUMERUS
C2853864|T191|C82.84|ICD10CM|OTHER TYPES OF FOLLICULAR LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB|OTH TYPES OF FOLICLAR LYMPH, NODES OF AXILLA AND UPPER LIMB
C2853865|T191|C82.85|ICD10CM|OTHER TYPES OF FOLLICULAR LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|OTH TYPES OF FOLICLAR LYMPH, NODES OF ING RGN AND LOWER LIMB
C2853866|T191|C82.86|ICD10CM|OTHER TYPES OF FOLLICULAR LYMPHOMA, INTRAPELVIC LYMPH NODES|OTHER TYPES OF FOLLICULAR LYMPHOMA, INTRAPELVIC LYMPH NODES
C2853867|T191|C82.87|ICD10CM|OTHER TYPES OF FOLLICULAR LYMPHOMA, SPLEEN|OTHER TYPES OF FOLLICULAR LYMPHOMA, SPLEEN
C2853860|T191|C82.80|ICD10CM|OTHER TYPES OF FOLLICULAR LYMPHOMA, UNSPECIFIED SITE|OTHER TYPES OF FOLLICULAR LYMPHOMA, UNSPECIFIED SITE
C2853861|T191|C82.81|ICD10CM|OTHER TYPES OF FOLLICULAR LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK|OTH TYPES OF FOLICLAR LYMPH, NODES OF HEAD, FACE, AND NECK
C2853862|T191|C82.82|ICD10CM|OTHER TYPES OF FOLLICULAR LYMPHOMA, INTRATHORACIC LYMPH NODES|OTH TYPES OF FOLLICULAR LYMPHOMA, INTRATHORACIC LYMPH NODES
C2853863|T191|C82.83|ICD10CM|OTHER TYPES OF FOLLICULAR LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES|OTH TYPES OF FOLLICULAR LYMPHOMA, INTRA-ABD LYMPH NODES
C2832682|T037|S06.9X2S|ICD10CM|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|UNSP INTRACRANIAL INJURY W LOC OF 31-59 MIN, SEQUELA
C2882947|T047|I70.641|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF THIGH|ATHSCL NONBIOL BYPASS OF THE LEFT LEG W ULCERATION OF THIGH
C2887301|T047|I87.312|ICD10CM|CHRONIC VENOUS HYPERTENSION (IDIOPATHIC) WITH ULCER OF LEFT LOWER EXTREMITY|CHRONIC VENOUS HYPERTENSION W ULCER OF L LOW EXTREM
C2887302|T047|I87.313|ICD10CM|CHRONIC VENOUS HYPERTENSION (IDIOPATHIC) WITH ULCER OF BILATERAL LOWER EXTREMITY|CHRONIC VENOUS HYPERTENSION W ULCER OF BILATERAL LOW EXTRM
C2853868|T191|C82.88|ICD10CM|OTHER TYPES OF FOLLICULAR LYMPHOMA, LYMPH NODES OF MULTIPLE SITES|OTH TYPES OF FOLLICULAR LYMPHOMA, LYMPH NODES MULT SITE
C2853869|T191|C82.89|ICD10CM|OTHER TYPES OF FOLLICULAR LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES|OTH TYPES OF FOLICLAR LYMPH, EXTRNOD AND SOLID ORGAN SITES
C2838387|T037|S32.512B|ICD10CM|FRACTURE OF SUPERIOR RIM OF LEFT PUBIS, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF SUPERIOR RIM OF LEFT PUBIS, INIT FOR OPN FX
C2832680|T037|S06.9X2A|ICD10CM|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|UNSP INTRACRANIAL INJURY W LOC OF 31-59 MIN, INIT
C2888847|T047|M00.159|ICD10CM|PNEUMOCOCCAL ARTHRITIS, UNSPECIFIED HIP|PNEUMOCOCCAL ARTHRITIS, UNSPECIFIED HIP
C2888846|T047|M00.152|ICD10CM|PNEUMOCOCCAL ARTHRITIS, LEFT HIP|PNEUMOCOCCAL ARTHRITIS, LEFT HIP
C2888845|T047|M00.151|ICD10CM|PNEUMOCOCCAL ARTHRITIS, RIGHT HIP|PNEUMOCOCCAL ARTHRITIS, RIGHT HIP
C2832222|T037|S06.340S|ICD10CM|TRAUMATIC HEMORRHAGE OF RIGHT CEREBRUM WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|TRAUM HEMOR RIGHT CEREBRUM W/O LOC, SEQUELA
C2832481|T037|S06.5X3A|ICD10CM|TRAUMATIC SUBDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|TRAUM SUBDR HEM W LOC OF 1-5 HRS 59 MIN, INIT
C3696797|T047|M08.88|ICD10CM|OTHER JUVENILE ARTHRITIS, OTHER SPECIFIED SITE|OTHER JUVENILE ARTHRITIS, OTHER SPECIFIED SITE
C0837740|T047|M08.89|ICD10AM|OTHER JUVENILE ARTHRITIS, MULTIPLE SITES|OTHER JUVENILE ARTHRITIS, SITE UNSPECIFIED
C0837740|T047||ICD10CM|OTHER JUVENILE ARTHRITIS, UNSPECIFIED SITE
C2832220|T037|S06.340A|ICD10CM|TRAUMATIC HEMORRHAGE OF RIGHT CEREBRUM WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|TRAUM HEMOR RIGHT CEREBRUM W/O LOSS OF CONSCIOUSNESS, INIT
C2832483|T037|S06.5X3S|ICD10CM|TRAUMATIC SUBDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, SEQUELA|TRAUM SUBDR HEM W LOC OF 1-5 HRS 59 MIN, SEQUELA
C2873852|T047|D86.84|ICD10CM|SARCOID PYELONEPHRITIS|SARCOID PYELONEPHRITIS
C0553718|T047|N28.0|ICD10CM|ISCHEMIA AND INFARCTION OF KIDNEY|RENAL ARTERY OCCLUSION
C0451646|T047|D86.82|ICD10CM|MULTIPLE CRANIAL NERVE PALSIES IN SARCOIDOSIS|MULTIPLE CRANIAL NERVE PALSIES IN SARCOIDOSIS
C2895204|T047|M35.04|ICD10CM|SICCA SYNDROME WITH TUBULO-INTERSTITIAL NEPHROPATHY|SICCA SYNDROME WITH TUBULO-INTERSTITIAL NEPHROPATHY
C0086981|T047|M35.00|ICD10CM|SICCA SYNDROME, UNSPECIFIED|SICCA SYNDROME, UNSPECIFIED
C2895200|T047|M35.01|ICD10CM|SICCA SYNDROME WITH KERATOCONJUNCTIVITIS|SICCA SYNDROME WITH KERATOCONJUNCTIVITIS
C2895201|T047|M35.02|ICD10CM|SICCA SYNDROME WITH LUNG INVOLVEMENT|SICCA SYNDROME WITH LUNG INVOLVEMENT
C2895202|T047|M35.03|ICD10CM|SICCA SYNDROME WITH MYOPATHY|SICCA SYNDROME WITH MYOPATHY
C2895205|T047|M35.09|ICD10CM|SICCA SYNDROME WITH OTHER ORGAN INVOLVEMENT|SICCA SYNDROME WITH OTHER ORGAN INVOLVEMENT
C2869891|T037|S98.912A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT FOOT, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF LEFT FOOT, LEVEL UNSP, INIT
C2888894|T047|M00.80|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, UNSPECIFIED JOINT|ARTHRITIS DUE TO OTHER BACTERIA, UNSPECIFIED JOINT
C2901842|T047|M86.312|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, LEFT SHOULDER|CHRONIC MULTIFOCAL OSTEOMYELITIS, LEFT SHOULDER
C2901841|T047|M86.311|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, RIGHT SHOULDER|CHRONIC MULTIFOCAL OSTEOMYELITIS, RIGHT SHOULDER
C2901922|T047|M86.641|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, RIGHT HAND|OTHER CHRONIC OSTEOMYELITIS, RIGHT HAND
C2901923|T047|M86.642|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, LEFT HAND|OTHER CHRONIC OSTEOMYELITIS, LEFT HAND
C2888925|T047|M00.88|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, VERTEBRAE|ARTHRITIS DUE TO OTHER BACTERIA, VERTEBRAE
C2888926|T047|M00.89|ICD10CM|POLYARTHRITIS DUE TO OTHER BACTERIA|POLYARTHRITIS DUE TO OTHER BACTERIA
C2901843|T047|M86.319|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, UNSPECIFIED SHOULDER|CHRONIC MULTIFOCAL OSTEOMYELITIS, UNSPECIFIED SHOULDER
C2901924|T047|M86.649|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, UNSPECIFIED HAND|OTHER CHRONIC OSTEOMYELITIS, UNSPECIFIED HAND
C2887934|T047|K72.10|ICD10CM|CHRONIC HEPATIC FAILURE WITHOUT COMA|CHRONIC HEPATIC FAILURE WITHOUT COMA
C1260406|T047|G31.09|ICD10CM|OTHER FRONTOTEMPORAL DEMENTIA|OTHER FRONTOTEMPORAL DEMENTIA
C1386519|T046||ICD10CM|PICK'S DISEASE
C2873943|T047|E08.649|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH HYPOGLYCEMIA WITHOUT COMA|DIABETES DUE TO UNDERLYING CONDITION W HYPOGLYCEMIA W/O COMA
C2891281|T037||ICD10CM|LIVER TRANSPLANT INFECTION
C2873942|T047|E08.641|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH HYPOGLYCEMIA WITH COMA|DIABETES DUE TO UNDERLYING CONDITION W HYPOGLYCEMIA W COMA
C1956097|T047|Q93.3|DMDICD10|DELETION OF SHORT ARM OF CHROMOSOME 4|DELETION DES KURZEN ARMES DES CHROMOSOMS 4
C2910368|T049|Q93.2|ICD10CM|CHROMOSOME REPLACED WITH RING, DICENTRIC OR ISOCHROMOSOME|CHROMOSOME REPLACED WITH RING, DICENTRIC OR ISOCHROMOSOME
C0432438|T047|Q93.1|DMDICD10|WHOLE CHROMOSOME MONOSOMY, MOSAICISM (MITOTIC NONDISJUNCTION)|VOLLSTAENDIGE MONOSOMIE, MOSAIK (MITOTISCHE NON-DISJUNCTION)
C2910367|T047|Q93.0|ICD10CM|WHOLE CHROMOSOME MONOSOMY, NONMOSAICISM (MEIOTIC NONDISJUNCTION)|WHOLE CHROMOSOME MONOSOMY,NONMOSAIC (MEIOTIC NONDISJUNCTION)
C1112486|T191||ICD10CM|AGGRESSIVE SYSTEMIC MASTOCYTOSIS
C4509018|T191|C96.20|ICD10CM|MALIGNANT MAST CELL NEOPLASM, UNSPECIFIED|MALIGNANT MAST CELL NEOPLASM, UNSPECIFIED
C2854107|T191|C91.51|ICD10CM|ADULT T-CELL LYMPHOMA/LEUKEMIA (HTLV-1-ASSOCIATED), IN REMISSION|ADULT T-CELL LYMPHOMA/LEUKEMIA (HTLV-1-ASSOC), IN REMISSION
C2854106|T191|C91.50|ICD10CM|ADULT T-CELL LYMPHOMA/LEUKEMIA (HTLV-1-ASSOCIATED) NOT HAVING ACHIEVED REMISSION|ADULT T-CELL LYMPH/LEUK (HTLV-1-ASSOC) NOT ACHIEVE REMISSION
C0495652|T049|Q93.9|DMDICD10|DELETION FROM AUTOSOMES, UNSPECIFIED|DELETION DER AUTOSOMEN, NICHT NAEHER BEZEICHNET
C2874044|T047|E10.39|ICD10CM|TYPE 1 DIABETES MELLITUS WITH OTHER DIABETIC OPHTHALMIC COMPLICATION|TYPE 1 DIABETES W OTH DIABETIC OPHTHALMIC COMPLICATION
C4480966|T191|C96.29|ICD10CM|OTHER MALIGNANT MAST CELL NEOPLASM|OTHER MALIGNANT MAST CELL NEOPLASM
C2833524|T037|S12.501A|ICD10CM|UNSPECIFIED NONDISPLACED FRACTURE OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP NONDISP FX OF SIXTH CERVICAL VERTEBRA, INIT FOR CLOS FX
C2832435|T037|S06.4X1S|ICD10CM|EPIDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|EPIDURAL HEMORRHAGE W LOC OF 30 MINUTES OR LESS, SEQUELA
C2833525|T037|S12.501B|ICD10CM|UNSPECIFIED NONDISPLACED FRACTURE OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP NONDISP FX OF SIXTH CERVICAL VERTEBRA, INIT FOR OPN FX
C2882419|T047|I65.03|ICD10CM|OCCLUSION AND STENOSIS OF BILATERAL VERTEBRAL ARTERIES|OCCLUSION AND STENOSIS OF BILATERAL VERTEBRAL ARTERIES
C2882307|T047|I60.50|ICD10CM|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM UNSPECIFIED VERTEBRAL ARTERY|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM UNSP VERTEB ART
C2882417|T047|I65.01|ICD10CM|OCCLUSION AND STENOSIS OF RIGHT VERTEBRAL ARTERY|OCCLUSION AND STENOSIS OF RIGHT VERTEBRAL ARTERY
C2882309|T047|I60.52|ICD10CM|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM LEFT VERTEBRAL ARTERY|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM L VERTEB ART
C2882420|T047|I65.09|ICD10CM|OCCLUSION AND STENOSIS OF UNSPECIFIED VERTEBRAL ARTERY|OCCLUSION AND STENOSIS OF UNSPECIFIED VERTEBRAL ARTERY
C2832433|T037|S06.4X1A|ICD10CM|EPIDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|EPIDURAL HEMORRHAGE W LOC OF 30 MINUTES OR LESS, INIT
C4269543|T037|S02.652S|ICD10CM|FRACTURE OF ANGLE OF LEFT MANDIBLE, SEQUELA|FRACTURE OF ANGLE OF LEFT MANDIBLE, SEQUELA
C2885191|T037|T61.8X2S|ICD10CM|TOXIC EFFECT OF OTHER SEAFOOD, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF OTH SEAFOOD, INTENTIONAL SELF-HARM, SEQUELA
C2884691|T037|T57.3X2S|ICD10CM|TOXIC EFFECT OF HYDROGEN CYANIDE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF HYDROGEN CYANIDE, SELF-HARM, SEQUELA
C2857105|T037|S72.101C|ICD10CM|UNSPECIFIED TROCHANTERIC FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP TROCHAN FX RIGHT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2857104|T037|S72.101B|ICD10CM|UNSPECIFIED TROCHANTERIC FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP TROCHAN FX RIGHT FEMUR, INIT FOR OPN FX TYPE I/2
C2857103|T037|S72.101A|ICD10CM|UNSPECIFIED TROCHANTERIC FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP TROCHANTERIC FRACTURE OF RIGHT FEMUR, INIT FOR CLOS FX
C2855902|T037|S68.119S|ICD10CM|COMPLETE TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF UNSPECIFIED FINGER, SEQUELA|COMPLETE TRAUMATIC MCP AMPUTATION OF UNSP FINGER, SEQUELA
C2891206|T037|T85.691S|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTRAPERITONEAL DIALYSIS CATHETER, SEQUELA|MECH COMPL OF INTRAPERITONEAL DIALYSIS CATHETER, SEQUELA
C2885189|T037|T61.8X2A|ICD10CM|TOXIC EFFECT OF OTHER SEAFOOD, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF OTH SEAFOOD, INTENTIONAL SELF-HARM, INIT
C2905655|T037|X71.2XXD|ICD10CM|INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION AFTER JUMP INTO SWIMMING POOL, SUBSEQUENT ENCOUNTER|SELF-HARM BY DROWN AFTER JUMP INTO SWIMMING POOL, SUBS
C2905654|T037|X71.2XXA|ICD10CM|INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION AFTER JUMP INTO SWIMMING POOL, INITIAL ENCOUNTER|SELF-HARM BY DROWN AFTER JUMP INTO SWIMMING POOL, INIT
C0268579|T047|E71.121|ICD10CM|PROPIONIC ACIDEMIA|PROPIONIC ACIDEMIA
C2869892|T037|S98.912D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT FOOT, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF LEFT FOOT, LEVEL UNSP, SUBS
C2905656|T037|X71.2XXS|ICD10CM|INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION AFTER JUMP INTO SWIMMING POOL, SEQUELA|SELF-HARM BY DROWN AFTER JUMP INTO SWIMMING POOL, SEQUELA
C0260762|T033|Z43.2|DMDICD10|ENCOUNTER FOR ATTENTION TO ILEOSTOMY|VERSORGUNG EINES ILEOSTOMAS
C2901205|T046|M84.534A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, LEFT RADIUS, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, LEFT RADIUS, INIT
C2887469|T047||ICD10CM|BRONCHIECTASIS, UNCOMPLICATED
C2896735|T046|M80.842A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, LEFT HAND, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, LEFT HAND, INIT
C2896720|T046|M80.839A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, UNSPECIFIED FOREARM, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, UNSP FOREARM, INIT
C2857259|T037|S72.121C|ICD10CM|DISPLACED FRACTURE OF LESSER TROCHANTER OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF LESS TROCHANTER OF R FEMR, 7THC
C2857258|T037|S72.121B|ICD10CM|DISPLACED FRACTURE OF LESSER TROCHANTER OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF LESS TROCHANTER OF R FEMR, 7THB
C0878696|T047||ICD10CM|BRONCHIECTASIS WITH (ACUTE) EXACERBATION
C2869856|T037|S98.229D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF TWO OR MORE UNSPECIFIED LESSER TOES, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMP OF TWO OR MORE UNSP LESSER TOES, SUBS
C2845900|T191|C69.01|ICD10CM|MALIGNANT NEOPLASM OF RIGHT CONJUNCTIVA|MALIGNANT NEOPLASM OF RIGHT CONJUNCTIVA
C2845899|T191|C69.00|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED CONJUNCTIVA|MALIGNANT NEOPLASM OF UNSPECIFIED CONJUNCTIVA
C2845901|T191|C69.02|ICD10CM|MALIGNANT NEOPLASM OF LEFT CONJUNCTIVA|MALIGNANT NEOPLASM OF LEFT CONJUNCTIVA
C2855947|T037|S68.411A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT HAND AT WRIST LEVEL, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMP OF RIGHT HAND AT WRIST LEVEL, INIT
C2877073|T037|T38.3X2S|ICD10CM|POISONING BY INSULIN AND ORAL HYPOGLYCEMIC [ANTIDIABETIC] DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY INSULIN AND ORAL HYPOGLYCEMIC DRUGS, SLF-HRM, SQLA
C2875341|T047|G82.53|ICD10CM|QUADRIPLEGIA, C5-C7 COMPLETE|QUADRIPLEGIA, C5-C7 COMPLETE
C2875340|T047|G82.52|ICD10CM|QUADRIPLEGIA, C1-C4 INCOMPLETE|QUADRIPLEGIA, C1-C4 INCOMPLETE
C2875339|T047|G82.51|ICD10CM|QUADRIPLEGIA, C1-C4 COMPLETE|QUADRIPLEGIA, C1-C4 COMPLETE
C0034372|T047|G82.5|ICD10AM|QUADRIPLEGIA, UNSPECIFIED|TETRAPLEGIA, UNSPECIFIED
C2875342|T047|G82.54|ICD10CM|QUADRIPLEGIA, C5-C7 INCOMPLETE|QUADRIPLEGIA, C5-C7 INCOMPLETE
C2889433|T047|M06.262|ICD10CM|RHEUMATOID BURSITIS, LEFT KNEE|RHEUMATOID BURSITIS, LEFT KNEE
C2889432|T047|M06.261|ICD10CM|RHEUMATOID BURSITIS, RIGHT KNEE|RHEUMATOID BURSITIS, RIGHT KNEE
C2901481|T046|M84.651A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, RIGHT FEMUR, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, RIGHT FEMUR, INIT
C2877071|T037|T38.3X2A|ICD10CM|POISONING BY INSULIN AND ORAL HYPOGLYCEMIC [ANTIDIABETIC] DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY INSULIN AND ORAL HYPOGLYCEMIC DRUGS, SLF-HRM, INIT
C2888945|T047|M01.X49|ICD10CM|DIRECT INFECTION OF UNSPECIFIED HAND IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIRECT INFCT OF UNSP HAND IN INFEC/PARASTC DIS CLASSD ELSWHR
C2889434|T047|M06.269|ICD10CM|RHEUMATOID BURSITIS, UNSPECIFIED KNEE|RHEUMATOID BURSITIS, UNSPECIFIED KNEE
C2888944|T047|M01.X42|ICD10CM|DIRECT INFECTION OF LEFT HAND IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIRECT INFCT OF L HAND IN INFEC/PARASTC DIS CLASSD ELSWHR
C2888943|T047|M01.X41|ICD10CM|DIRECT INFECTION OF RIGHT HAND IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIRECT INFCT OF R HAND IN INFEC/PARASTC DIS CLASSD ELSWHR
C4269419|T037|S02.600A|ICD10CM|FRACTURE OF UNSPECIFIED PART OF BODY OF MANDIBLE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FX UNSP PART OF BODY OF MANDIBLE, UNSPECIFIED SIDE, INIT
C2890342|T037|T83.420A|ICD10CM|DISPLACEMENT OF IMPLANTED PENILE PROSTHESIS, INITIAL ENCOUNTER|DISPLACEMENT OF IMPLANTED PENILE PROSTHESIS, INIT
C2837775|T037|S32.16XB|ICD10CM|TYPE 3 FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE 3 FRACTURE OF SACRUM, INIT ENCNTR FOR OPEN FRACTURE
C2837774|T037|S32.16XA|ICD10CM|TYPE 3 FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE 3 FRACTURE OF SACRUM, INIT ENCNTR FOR CLOSED FRACTURE
C0838504|T047|M46.22|ICD10AM|OSTEOMYELITIS OF VERTEBRA, CERVICAL REGION|OSTEOMYELITIS OF VERTEBRA, CERVICAL REGION
C0838505|T047|M46.23|ICD10AM|OSTEOMYELITIS OF VERTEBRA, CERVICOTHORACIC REGION|OSTEOMYELITIS OF VERTEBRA, CERVICOTHORACIC REGION
C2883586|T037|T50.2X2S|ICD10CM|POISONING BY CARBONIC-ANHYDRASE INHIBITORS, BENZOTHIADIAZIDES AND OTHER DIURETICS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY CRBNC-ANHYDR INHIBTR,BENZO/OTH DIURETC,SLF-HRM,SQLA
C0838506|T047|M46.24|ICD10AM|OSTEOMYELITIS OF VERTEBRA, THORACIC REGION|OSTEOMYELITIS OF VERTEBRA, THORACIC REGION
C2883334|T037|T49.2X2S|ICD10CM|POISONING BY LOCAL ASTRINGENTS AND LOCAL DETERGENTS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY LOCAL ASTRINGENTS/DETERGENTS, SELF-HARM, SEQUELA
C2242796|T047|D57.40|ICD10CM|SICKLE-CELL THALASSEMIA WITHOUT CRISIS|MICRODREPANOCYTOSIS
C2883332|T037|T49.2X2A|ICD10CM|POISONING BY LOCAL ASTRINGENTS AND LOCAL DETERGENTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY LOCAL ASTRINGENTS/DETERGENTS, SELF-HARM, INIT
C0153413|T191|C15.3|DMDICD10|MALIGNANT NEOPLASM OF UPPER THIRD OF ESOPHAGUS|BOESARTIGE NEUBILDUNG: OESOPHAGUS, OBERES DRITTEL
C0153415|T191|C15.5|DMDICD10|MALIGNANT NEOPLASM OF LOWER THIRD OF ESOPHAGUS|BOESARTIGE NEUBILDUNG: OESOPHAGUS, UNTERES DRITTEL
C0153414|T191|C15.4|DMDICD10|MALIGNANT NEOPLASM OF MIDDLE THIRD OF ESOPHAGUS|BOESARTIGE NEUBILDUNG: OESOPHAGUS, MITTLERES DRITTEL
C2901169|T046|M84.522A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, LEFT HUMERUS, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, L HUMERUS, INIT
C2905684|T037|X73.2XXD|ICD10CM|INTENTIONAL SELF-HARM BY MACHINE GUN DISCHARGE, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY MACHINE GUN DISCHARGE, SUBS ENCNTR
C0546837|T191|C15.9|DMDICD10|MALIGNANT NEOPLASM OF ESOPHAGUS, UNSPECIFIED|BOESARTIGE NEUBILDUNG: OESOPHAGUS, NICHT NAEHER BEZEICHNET
C0496776|T191|C15.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF ESOPHAGUS|BOESARTIGE NEUBILDUNG: OESOPHAGUS, MEHRERE TEILBEREICHE UEBERLAPPEND
C2832383|T037|S06.379A|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF CEREBELLUM WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|CONTUS/LAC/HEM CRBLM W LOC OF UNSP DURATION, INIT
C2902038|T046|M87.221|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, RIGHT HUMERUS|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, RIGHT HUMERUS
C2888643|T047|L97.109|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED THIGH WITH UNSPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF UNSP THIGH WITH UNSP SEVERITY
C4509277|T047|L97.108|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED THIGH WITH OTHER SPECIFIED SEVERITY|NON-PRS CHRONIC ULCER OF UNSPECIFIED THIGH WITH OTH SEVERITY
C4509276|T047|L97.106|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED THIGH WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OF UNSP THIGH WITH BONE INVL W/O EVD OF NECR
C4509275|T047|L97.105|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED THIGH WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OF UNSP THIGH WITH MSL INVL W/O EVD OF NECR
C2888642|T047|L97.104|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED THIGH WITH NECROSIS OF BONE|NON-PRESSURE CHRONIC ULCER OF UNSP THIGH W NECROSIS OF BONE
C2888641|T047|L97.103|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED THIGH WITH NECROSIS OF MUSCLE|NON-PRS CHRONIC ULCER OF UNSP THIGH W NECROSIS OF MUSCLE
C2888640|T047|L97.102|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED THIGH WITH FAT LAYER EXPOSED|NON-PRESSURE CHRONIC ULCER OF UNSP THIGH W FAT LAYER EXPOSED
C2888639|T047|L97.101|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED THIGH LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHRONIC ULCER OF UNSP THIGH LIMITED TO BRKDWN SKIN
C2977869|T037|S32.592A|ICD10CM|OTHER SPECIFIED FRACTURE OF LEFT PUBIS, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF LEFT PUBIS, INIT ENCNTR FOR CLOSED FRACTURE
C2902925|T047|N07.9|ICD10CM|HEREDITARY NEPHROPATHY, NOT ELSEWHERE CLASSIFIED WITH UNSPECIFIED MORPHOLOGIC LESIONS|HEREDITARY NEPHROPATHY, NEC W UNSP MORPHOLOGIC LESIONS
C2902924|T047|N07.8|ICD10CM|HEREDITARY NEPHROPATHY, NOT ELSEWHERE CLASSIFIED WITH OTHER MORPHOLOGIC LESIONS|HEREDITARY NEPHROPATHY, NEC W OTH MORPHOLOGIC LESIONS
C2902922|T047|N07.7|ICD10CM|HEREDITARY NEPHROPATHY, NOT ELSEWHERE CLASSIFIED WITH DIFFUSE CRESCENTIC GLOMERULONEPHRITIS|HEREDITARY NEPHROPATHY, NOT ELSEWHERE CLASSIFIED WITH EXTRACAPILLARY GLOMERULONEPHRITIS
C2902921|T047|N07.6|ICD10CM|HEREDITARY NEPHROPATHY, NOT ELSEWHERE CLASSIFIED WITH DENSE DEPOSIT DISEASE|HEREDITARY NEPHROPATHY, NOT ELSEWHERE CLASSIFIED WITH MEMBRANOPROLIFERATIVE GLOMERULONEPHRITIS, TYPE 2
C2902920|T047|N07.5|ICD10CM|HEREDITARY NEPHROPATHY, NOT ELSEWHERE CLASSIFIED WITH DIFFUSE MESANGIOCAPILLARY GLOMERULONEPHRITIS|HEREDITARY NEPHROPATHY, NOT ELSEWHERE CLASSIFIED WITH MEMBRANOPROLIFERATIVE GLOMERULONEPHRITIS, TYPES 1 AND 3, OR NOS
C0868880|T047|N07.4|DMDICD10|HEREDITARY NEPHROPATHY, NOT ELSEWHERE CLASSIFIED WITH DIFFUSE ENDOCAPILLARY PROLIFERATIVE GLOMERULONEPHRITIS|HEREDITAERE NEPHROPATHIE, ANDERENORTS NICHT KLASSIFIZIERT: DIFFUSE ENDOKAPILLAER-PROLIFERATIVE GLOMERULONEPHRITIS
C0868878|T047|N07.3|DMDICD10|HEREDITARY NEPHROPATHY, NOT ELSEWHERE CLASSIFIED WITH DIFFUSE MESANGIAL PROLIFERATIVE GLOMERULONEPHRITIS|HEREDITAERE NEPHROPATHIE, ANDERENORTS NICHT KLASSIFIZIERT: DIFFUSE MESANGIOPROLIFERATIVE GLOMERULONEPHRITIS
C0868875|T047|N07.2|DMDICD10|HEREDITARY NEPHROPATHY, NOT ELSEWHERE CLASSIFIED WITH DIFFUSE MEMBRANOUS GLOMERULONEPHRITIS|HEREDITAERE NEPHROPATHIE, ANDERENORTS NICHT KLASSIFIZIERT: DIFFUSE MEMBRANOESE GLOMERULONEPHRITIS
C2902919|T047|N07.1|ICD10CM|HEREDITARY NEPHROPATHY, NOT ELSEWHERE CLASSIFIED WITH FOCAL AND SEGMENTAL GLOMERULAR LESIONS|HEREDITARY NEPHROPATHY, NOT ELSEWHERE CLASSIFIED WITH FOCAL GLOMERULONEPHRITIS
C2902916|T047|N07.0|ICD10CM|HEREDITARY NEPHROPATHY, NOT ELSEWHERE CLASSIFIED WITH MINOR GLOMERULAR ABNORMALITY|HEREDITARY NEPHROPATHY, NOT ELSEWHERE CLASSIFIED WITH MINIMAL CHANGE LESION
C2890883|T037|T84.629A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL FIXATION DEVICE OF UNSPECIFIED BONE OF LEG, INITIAL ENCOUNTER|INFECT/INFLM REACT DUE TO INT FIX OF UNSP BONE OF LEG, INIT
C0153754|T191|C81.43|ICD10CM|LYMPHOCYTE-RICH HODGKIN LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES|LYMPHOCYTE-RICH HODGKIN LYMPHOMA, INTRA-ABD LYMPH NODES
C0153753|T191||ICD10CM|LYMPHOCYTE-RICH HODGKIN LYMPHOMA, INTRATHORACIC LYMPH NODES
C4267863|T191|C81.41|ICD10CM|LYMPHOCYTE-RICH HODGKIN LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK|LYMP-RICH HODGKIN LYMPHOMA, NODES OF HEAD, FACE, AND NECK
C4267862|T191|C81.40|ICD10CM|LYMPHOCYTE-RICH HODGKIN LYMPHOMA, UNSPECIFIED SITE|LYMPHOCYTE-RICH HODGKIN LYMPHOMA, UNSPECIFIED SITE
C0153758|T191||ICD10CM|LYMPHOCYTE-RICH HODGKIN LYMPHOMA, SPLEEN
C0153757|T191||ICD10CM|LYMPHOCYTE-RICH HODGKIN LYMPHOMA, INTRAPELVIC LYMPH NODES
C4267865|T191|C81.45|ICD10CM|LYMPHOCYTE-RICH HODGKIN LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|LYMP-RICH HODGKIN LYMPH, NODES OF ING REGION AND LOWER LIMB
C4267864|T191|C81.44|ICD10CM|LYMPHOCYTE-RICH HODGKIN LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB|LYMP-RICH HODGKIN LYMPHOMA, NODES OF AXILLA AND UPPER LIMB
C2838258|T037|S32.466B|ICD10CM|NONDISPLACED ASSOCIATED TRANSVERSE-POSTERIOR FRACTURE OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP ASSOC TRANSV/POST FX UNSP ACETAB, INIT FOR OPN FX
C4267866|T191|C81.49|ICD10CM|LYMPHOCYTE-RICH HODGKIN LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES|LYMP-RICH HODGKIN LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES
C0153759|T191|C81.48|ICD10CM|LYMPHOCYTE-RICH HODGKIN LYMPHOMA, LYMPH NODES OF MULTIPLE SITES|LYMPHOCYTE-RICH HODGKIN LYMPHOMA, LYMPH NODES MULT SITE
C4268219|T048|F12.288|ICD10CM|CANNABIS DEPENDENCE WITH OTHER CANNABIS-INDUCED DISORDER|CANNABIS USE DISORDER, SEVERE, WITH CANNABIS-INDUCED SLEEP DISORDER
C2889018|T047|M02.172|ICD10CM|POSTDYSENTERIC ARTHROPATHY, LEFT ANKLE AND FOOT|POSTDYSENTERIC ARTHROPATHY, LEFT ANKLE AND FOOT
C2889017|T047|M02.171|ICD10CM|POSTDYSENTERIC ARTHROPATHY, RIGHT ANKLE AND FOOT|POSTDYSENTERIC ARTHROPATHY, RIGHT ANKLE AND FOOT
C2833949|T037|S14.128S|ICD10CM|CENTRAL CORD SYNDROME AT C8 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|CENTRAL CORD SYNDROME AT C8, SEQUELA
C2889019|T047|M02.179|ICD10CM|POSTDYSENTERIC ARTHROPATHY, UNSPECIFIED ANKLE AND FOOT|POSTDYSENTERIC ARTHROPATHY, UNSPECIFIED ANKLE AND FOOT
C0340530|T046|T86.21|ICD10CM|HEART TRANSPLANT REJECTION|HEART TRANSPLANT REJECTION
C2891272|T037|T86.20|ICD10CM|UNSPECIFIED COMPLICATION OF HEART TRANSPLANT|UNSPECIFIED COMPLICATION OF HEART TRANSPLANT
C2891273|T037||ICD10CM|HEART TRANSPLANT INFECTION
C0340531|T046||ICD10CM|HEART TRANSPLANT FAILURE
C2884432|T037|T55.0X2S|ICD10CM|TOXIC EFFECT OF SOAPS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF SOAPS, INTENTIONAL SELF-HARM, SEQUELA
C2891280|T037|T86.40|ICD10CM|UNSPECIFIED COMPLICATION OF LIVER TRANSPLANT|UNSPECIFIED COMPLICATION OF LIVER TRANSPLANT
C2879772|T037|T47.4X2A|ICD10CM|POISONING BY OTHER LAXATIVES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH LAXATIVES, INTENTIONAL SELF-HARM, INIT
C2838042|T037|S32.416A|ICD10CM|NONDISPLACED FRACTURE OF ANTERIOR WALL OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF ANTERIOR WALL OF UNSP ACETABULUM, INIT
C2837847|T037|S32.314B|ICD10CM|NONDISPLACED AVULSION FRACTURE OF RIGHT ILIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP AVULSION FRACTURE OF RIGHT ILIUM, INIT FOR OPN FX
C2837846|T037|S32.314A|ICD10CM|NONDISPLACED AVULSION FRACTURE OF RIGHT ILIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED AVULSION FRACTURE OF RIGHT ILIUM, INIT
C2884430|T037|T55.0X2A|ICD10CM|TOXIC EFFECT OF SOAPS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF SOAPS, INTENTIONAL SELF-HARM, INIT ENCNTR
C2838365|T037|S32.499A|ICD10CM|OTHER SPECIFIED FRACTURE OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF UNSP ACETABULUM, INIT FOR CLOS FX
C2888851|T047|M00.169|ICD10CM|PNEUMOCOCCAL ARTHRITIS, UNSPECIFIED KNEE|PNEUMOCOCCAL ARTHRITIS, UNSPECIFIED KNEE
C2977698|T037|S02.42XA|ICD10CM|FRACTURE OF ALVEOLUS OF MAXILLA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF ALVEOLUS OF MAXILLA, INIT FOR CLOS FX
C2977699|T037|S02.42XB|ICD10CM|FRACTURE OF ALVEOLUS OF MAXILLA, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF ALVEOLUS OF MAXILLA, INIT FOR OPN FX
C2874372|T048||ICD10CM|ALCOHOL ABUSE WITH INTOXICATION, UNCOMPLICATED
C2838157|T037|S32.444A|ICD10CM|NONDISPLACED FRACTURE OF POSTERIOR COLUMN [ILIOISCHIAL] OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF POSTERIOR COLUMN OF RIGHT ACETABULUM, INIT
C2837538|T037|S32.028A|ICD10CM|OTHER FRACTURE OF SECOND LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF SECOND LUMBAR VERTEBRA, INIT FOR CLOS FX
C2837539|T037|S32.028B|ICD10CM|OTHER FRACTURE OF SECOND LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF SECOND LUMBAR VERTEBRA, INIT FOR OPN FX
C2887155|T047|I82.B23|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF SUBCLAVIAN VEIN, BILATERAL|CHRONIC EMBOLISM AND THROMBOSIS OF SUBCLAV VEIN, BILATERAL
C2887154|T047|I82.B22|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF LEFT SUBCLAVIAN VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF LEFT SUBCLAVIAN VEIN
C2887153|T047|I82.B21|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF RIGHT SUBCLAVIAN VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF RIGHT SUBCLAVIAN VEIN
C2977703|T037|S02.42XS|ICD10CM|FRACTURE OF ALVEOLUS OF MAXILLA, SEQUELA|FRACTURE OF ALVEOLUS OF MAXILLA, SEQUELA
C2887156|T047|I82.B29|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED SUBCLAVIAN VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF UNSP SUBCLAVIAN VEIN
C2879774|T037|T47.4X2S|ICD10CM|POISONING BY OTHER LAXATIVES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTHER LAXATIVES, INTENTIONAL SELF-HARM, SEQUELA
C2873892|T047|E08.22|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH DIABETIC CHRONIC KIDNEY DISEASE|DIABETES DUE TO UNDRL COND W DIABETIC CHRONIC KIDNEY DISEASE
C2875189|T047|G43.919|ICD10CM|MIGRAINE, UNSPECIFIED, INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|MIGRAINE, UNSP, INTRACTABLE, WITHOUT STATUS MIGRAINOSUS
C2834032|T037|S14.151A|ICD10CM|OTHER INCOMPLETE LESION AT C1 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|OTH INCOMPLETE LESION AT C1, INIT
C2905650|T037|X71.1XXA|ICD10CM|INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION WHILE IN SWIMMING POOL, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY DROWN WHILE IN SWIMMING POOL, INIT
C2875188|T047|G43.911|ICD10CM|MIGRAINE, UNSPECIFIED, INTRACTABLE, WITH STATUS MIGRAINOSUS|MIGRAINE, UNSPECIFIED, INTRACTABLE, WITH STATUS MIGRAINOSUS
C2876695|T037|T36.6X2S|ICD10CM|POISONING BY RIFAMPICINS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY RIFAMPICINS, INTENTIONAL SELF-HARM, SEQUELA
C2886919|T037|T81.512A|ICD10CM|ADHESIONS DUE TO FOREIGN BODY ACCIDENTALLY LEFT IN BODY FOLLOWING KIDNEY DIALYSIS, INITIAL ENCOUNTER|ADHES DUE TO FB ACC LEFT IN BODY FOL KIDNEY DIALYSIS, INIT
C0864871|T191||ICD10CM|MALIGNANT NEOPLASM OF CECUM
C2874463|T048|F11.951|ICD10CM|OPIOID USE, UNSPECIFIED WITH OPIOID-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|OPIOID USE, UNSP W OPIOID-INDUC PSYCH DISORDER W HALLUCIN
C0153439|T191|C18.2|DMDICD10|MALIGNANT NEOPLASM OF ASCENDING COLON|BOESARTIGE NEUBILDUNG: COLON ASCENDENS
C0338952|T048|F48.1|DMDICD10|DEPERSONALIZATION-DEREALIZATION SYNDROME|DEPERSONALISATIONS- UND DEREALISATIONSSYNDROM
C2882513|T047|I69.163|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING RIGHT NON-DOMINANT SIDE|OTH PARLYT SYND FOL NTRM INTCRBL HEMOR AFF RIGHT NONDOM SIDE
C2882512|T047|I69.162|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING LEFT DOMINANT SIDE|OTH PARLYT SYNDROME FOL NTRM INTCRBL HEMOR AFF LEFT DOM SIDE
C2882511|T047|I69.161|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING RIGHT DOMINANT SIDE|OTH PARLYT SYND FOL NTRM INTCRBL HEMOR AFF RIGHT DOM SIDE
C2873871|T047|E05.30|ICD10CM|THYROTOXICOSIS FROM ECTOPIC THYROID TISSUE WITHOUT THYROTOXIC CRISIS OR STORM|THYROTXCOSIS FROM ECTOPIC THYROID TISSUE W/O THYROTXC CRISIS
C4237282|T048|F19.959|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH PSYCHOACTIVE SUBSTANCE-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|OTHER OR UNKNOWN SUBSTANCE-INDUCED PSYCHOTIC DISORDER, WITHOUT USE DISORDER
C2882515|T047|I69.165|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE, BILATERAL|OTH PARALYTIC SYNDROME FOLLOWING NTRM INTCRBL HEMOR, BI
C2882514|T047|I69.164|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING LEFT NON-DOMINANT SIDE|OTH PARLYT SYND FOL NTRM INTCRBL HEMOR AFF LEFT NONDOM SIDE
C2882362|T047|I63.30|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF UNSPECIFIED CEREBRAL ARTERY|CEREBRAL INFARCTION DUE TO THOMBOS UNSP CEREBRAL ARTERY
C2882516|T047|I69.169|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING UNSPECIFIED SIDE|OTH PARALYTIC SYNDROME FOL NTRM INTCRBL HEMOR AFF UNSP SIDE
C2874847|T048|F19.950|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH PSYCHOACTIVE SUBSTANCE-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|OTH PSYCHOACTV SUB USE, UNSP W PSYCH DISORDER W DELUSIONS
C2889484|T047|M06.859|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, UNSPECIFIED HIP|OTHER SPECIFIED RHEUMATOID ARTHRITIS, UNSPECIFIED HIP
C0431321|T019|Q05.0|DMDICD10|CERVICAL SPINA BIFIDA WITH HYDROCEPHALUS|ZERVIKALE SPINA BIFIDA MIT HYDROZEPHALUS
C1409928|T019||ICD10CM|THORACIC SPINA BIFIDA WITH HYDROCEPHALUS
C1409927|T019||ICD10CM|LUMBAR SPINA BIFIDA WITH HYDROCEPHALUS
C0495474|T019|Q05.3|DMDICD10|SACRAL SPINA BIFIDA WITH HYDROCEPHALUS|SAKRALE SPINA BIFIDA MIT HYDROZEPHALUS
C0477973|T019|Q05.4|DMDICD10|UNSPECIFIED SPINA BIFIDA WITH HYDROCEPHALUS|NICHT NAEHER BEZEICHNETE SPINA BIFIDA MIT HYDROZEPHALUS
C0158535|T019|Q05.5|DMDICD10|CERVICAL SPINA BIFIDA WITHOUT HYDROCEPHALUS|ZERVIKALE SPINA BIFIDA OHNE HYDROZEPHALUS
C1406918|T019||ICD10CM|THORACIC SPINA BIFIDA WITHOUT HYDROCEPHALUS
C1403241|T019||ICD10CM|LUMBAR SPINA BIFIDA WITHOUT HYDROCEPHALUS
C0495478|T019|Q05.8|DMDICD10|SACRAL SPINA BIFIDA WITHOUT HYDROCEPHALUS|SAKRALE SPINA BIFIDA OHNE HYDROZEPHALUS
C0080178|T019|Q05.9|DMDICD10|SPINA BIFIDA, UNSPECIFIED|SPINA BIFIDA, NICHT NAEHER BEZEICHNET
C2869807|T037|S98.131A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF ONE RIGHT LESSER TOE, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF ONE RIGHT LESSER TOE, INIT
C4290172|T047|I70.65|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF OTHER EXTREMITY WITH ULCERATION|ANY CONDITION CLASSIFIABLE TO I70.618 AND I70.628
C0346629|T191||ICD10CM|MALIGNANT NEOPLASM OF COLON, UNSPECIFIED
C0036980|T046|R57.0|DMDICD10|CARDIOGENIC SHOCK|KARDIOGENER SCHOCK
C0020683|T046|R57.1|DMDICD10|HYPOVOLEMIC SHOCK|HYPOVOLAEMISCHER SCHOCK
C4269300|T037|S02.11DA|ICD10CM|TYPE II OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE II OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, INIT
C4269301|T037|S02.11DB|ICD10CM|TYPE II OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE II OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, 7THB
C2869809|T037|S98.131S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF ONE RIGHT LESSER TOE, SEQUELA|COMPLETE TRAUMATIC AMP OF ONE RIGHT LESSER TOE, SEQUELA
C2832051|T037|S06.2X9S|ICD10CM|DIFFUSE TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|DIFFUSE TBI W LOC OF UNSP DURATION, SEQUELA
C2832426|T037|S06.389S|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF BRAINSTEM WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|CONTUS/LAC/HEM BRAINSTEM W LOC OF UNSP DURATION, SEQUELA
C2832113|T037|S06.314S|ICD10CM|CONTUSION AND LACERATION OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|CONTUS/LAC RIGHT CEREBRUM W LOC OF 6-24 HRS, SEQUELA
C2833458|T037|S12.401B|ICD10CM|UNSPECIFIED NONDISPLACED FRACTURE OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP NONDISP FX OF FIFTH CERVICAL VERTEBRA, INIT FOR OPN FX
C2830246|T047|B48.8|ICD10CM|OTHER SPECIFIED MYCOSES|INFECTION OF TISSUE AND ORGANS BY SAPROPHYTIC FUNGI NEC
C2833457|T037|S12.401A|ICD10CM|UNSPECIFIED NONDISPLACED FRACTURE OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP NONDISP FX OF FIFTH CERVICAL VERTEBRA, INIT FOR CLOS FX
C2832424|T037|S06.389A|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF BRAINSTEM WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|CONTUS/LAC/HEM BRAINSTEM W LOC OF UNSP DURATION, INIT
C0348993|T047|B48.4|DMDICD10|PENICILLOSIS|PENIZILLIOSE
C2869857|T037|S98.229S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF TWO OR MORE UNSPECIFIED LESSER TOES, SEQUELA|PARTIAL TRAUM AMP OF TWO OR MORE UNSP LESSER TOES, SEQUELA
C2902378|T047|M89.669|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, UNSPECIFIED LOWER LEG|OSTEOPATHY AFTER POLIOMYELITIS, UNSPECIFIED LOWER LEG
C2838115|T037|S32.434B|ICD10CM|NONDISPLACED FRACTURE OF ANTERIOR COLUMN [ILIOPUBIC] OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP FX OF ANT COLUMN OF RIGHT ACETAB, INIT FOR OPN FX
C2887781|T047|K50.911|ICD10CM|CROHN'S DISEASE, UNSPECIFIED, WITH RECTAL BLEEDING|CROHN'S DISEASE, UNSPECIFIED, WITH RECTAL BLEEDING
C2874173|T047|E13.638|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH OTHER ORAL COMPLICATIONS|OTH DIABETES MELLITUS WITH OTHER ORAL COMPLICATIONS
C2902377|T047|M89.662|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, LEFT LOWER LEG|OSTEOPATHY AFTER POLIOMYELITIS, LEFT LOWER LEG
C2874172|T047|E13.630|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PERIODONTAL DISEASE|OTHER SPECIFIED DIABETES MELLITUS WITH PERIODONTAL DISEASE
C2890213|T037|T83.020A|ICD10CM|DISPLACEMENT OF CYSTOSTOMY CATHETER, INITIAL ENCOUNTER|DISPLACEMENT OF CYSTOSTOMY CATHETER, INITIAL ENCOUNTER
C2902376|T047|M89.661|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, RIGHT LOWER LEG|OSTEOPATHY AFTER POLIOMYELITIS, RIGHT LOWER LEG
C2884915|T037|T59.5X2S|ICD10CM|TOXIC EFFECT OF FLUORINE GAS AND HYDROGEN FLUORIDE, INTENTIONAL SELF-HARM, SEQUELA|TOX EFF OF FLUORINE GAS AND HYDROGEN FLUORIDE, SLF-HRM, SQLA
C1400398|T020||ICD10CM|OTHER INTESTINAL OBSTRUCTION
C0021843|T047|K56.69|ICD10CM|UNSPECIFIED INTESTINAL OBSTRUCTION|OCCLUSION OF COLON OR INTESTINE NOS
C2887786|T047|K50.919|ICD10CM|CROHN'S DISEASE, UNSPECIFIED, WITH UNSPECIFIED COMPLICATIONS|CROHN'S DISEASE, UNSPECIFIED, WITH UNSPECIFIED COMPLICATIONS
C2902734|T037|M96.639|ICD10CM|FRACTURE OF RADIUS OR ULNA FOLLOWING INSERTION OF ORTHOPEDIC IMPLANT, JOINT PROSTHESIS, OR BONE PLATE, UNSPECIFIED ARM|FX RAD/ULNA FOL INSRT ORTHO IMPLNT/PROSTH/BONE PLT, UNSP ARM
C2889165|T047|M05.20|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE
C2902732|T037|M96.631|ICD10CM|FRACTURE OF RADIUS OR ULNA FOLLOWING INSERTION OF ORTHOPEDIC IMPLANT, JOINT PROSTHESIS, OR BONE PLATE, RIGHT ARM|FX RAD/ULNA FOL INSRT ORTHO IMPLNT/PROSTH/BONE PLT, R ARM
C2889195|T047|M05.29|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS MULT SITE
C2902733|T037|M96.632|ICD10CM|FRACTURE OF RADIUS OR ULNA FOLLOWING INSERTION OF ORTHOPEDIC IMPLANT, JOINT PROSTHESIS, OR BONE PLATE, LEFT ARM|FX RAD/ULNA FOL INSRT ORTHO IMPLNT/PROSTH/BONE PLT, LEFT ARM
C2901966|T046|M87.059|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED FEMUR|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED FEMUR
C2856499|T037|S72.002A|ICD10CM|FRACTURE OF UNSPECIFIED PART OF NECK OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF UNSP PART OF NECK OF LEFT FEMUR, INIT
C2901964|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF LEFT FEMUR
C2901963|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF RIGHT FEMUR
C2901962|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF PELVIS
C2886747|T037|T79.9XXA|ICD10CM|UNSPECIFIED EARLY COMPLICATION OF TRAUMA, INITIAL ENCOUNTER|UNSPECIFIED EARLY COMPLICATION OF TRAUMA, INITIAL ENCOUNTER
C2889350|T047|M05.769|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED KNEE WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRITIS W RHEU FACTOR OF UNSP KNEE W/O ORG/SYS INVOLV
C2889349|T047|M05.762|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT KNEE WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRITIS W RHEU FACTOR OF LEFT KNEE W/O ORG/SYS INVOLV
C2889348|T047|M05.761|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT KNEE WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRITIS W RHEU FACTOR OF R KNEE W/O ORG/SYS INVOLV
C2901242|T046|M84.550A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, PELVIS, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, PELVIS, INIT
C2887752|T047|K50.00|ICD10CM|CROHN'S DISEASE OF SMALL INTESTINE WITHOUT COMPLICATIONS|CROHN'S DISEASE OF SMALL INTESTINE WITHOUT COMPLICATIONS
C2882395|T047|I63.442|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF LEFT CEREBELLAR ARTERY|CEREBRAL INFARCTION DUE TO EMBOLISM OF LEFT CEREBLR ARTERY
C4268488|T047|I63.443|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF BILATERAL CEREBELLAR ARTERIES|CEREBRAL INFRC DUE TO EMBOLISM OF BILATERAL CEREBLR ARTERIES
C2882394|T047|I63.441|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF RIGHT CEREBELLAR ARTERY|CEREBRAL INFARCTION DUE TO EMBOLISM OF RIGHT CEREBLR ARTERY
C2882396|T047|I63.449|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF UNSPECIFIED CEREBELLAR ARTERY|CEREBRAL INFARCTION DUE TO EMBOLISM OF UNSP CEREBLR ARTERY
C2884705|T037|T57.8X2A|ICD10CM|TOXIC EFFECT OF OTHER SPECIFIED INORGANIC SUBSTANCES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF INORGANIC SUBSTANCES, SELF-HARM, INIT
C2875145|T047|G43.001|ICD10CM|MIGRAINE WITHOUT AURA, NOT INTRACTABLE, WITH STATUS MIGRAINOSUS|MIGRAINE W/O AURA, NOT INTRACTABLE, WITH STATUS MIGRAINOSUS
C2878020|T037|T41.5X2A|ICD10CM|POISONING BY THERAPEUTIC GASES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY THERAPEUTIC GASES, INTENTIONAL SELF-HARM, INIT
C2885919|T037|T63.892S|ICD10CM|TOXIC EFFECT OF CONTACT WITH OTHER VENOMOUS ANIMALS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CNTCT W OTH VENOM ANIMALS, SLF-HRM, SEQUELA
C2875146|T047|G43.009|ICD10CM|MIGRAINE WITHOUT AURA, NOT INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|MIGRAINE W/O AURA, NOT INTRACTABLE, W/O STATUS MIGRAINOSUS
C1955786|T046|I76|ICD10CM|SEPTIC ARTERIAL EMBOLISM|SEPTIC ARTERIAL EMBOLISM
C2884707|T037|T57.8X2S|ICD10CM|TOXIC EFFECT OF OTHER SPECIFIED INORGANIC SUBSTANCES, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF INORGANIC SUBSTANCES, SELF-HARM, SEQUELA
C2878022|T037|T41.5X2S|ICD10CM|POISONING BY THERAPEUTIC GASES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY THERAPEUTIC GASES, SELF-HARM, SEQUELA
C2885917|T037|T63.892A|ICD10CM|TOXIC EFFECT OF CONTACT WITH OTHER VENOMOUS ANIMALS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CONTACT W OTH VENOM ANIMALS, SLF-HRM, INIT
C2883433|T037|T49.6X2S|ICD10CM|POISONING BY OTORHINOLARYNGOLOGICAL DRUGS AND PREPARATIONS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTORHINO DRUGS AND PREP, SELF-HARM, SEQUELA
C2834046|T037|S14.154S|ICD10CM|OTHER INCOMPLETE LESION AT C4 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|OTH INCOMPLETE LESION AT C4, SEQUELA
C2883431|T037|T49.6X2A|ICD10CM|POISONING BY OTORHINOLARYNGOLOGICAL DRUGS AND PREPARATIONS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTORHINO DRUGS AND PREP, SELF-HARM, INIT
C4270266|T046|T83.123A|ICD10CM|DISPLACEMENT OF OTHER URINARY STENTS, INITIAL ENCOUNTER|DISPLACEMENT OF OTHER URINARY STENTS, INITIAL ENCOUNTER
C2834044|T037|S14.154A|ICD10CM|OTHER INCOMPLETE LESION AT C4 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|OTH INCOMPLETE LESION AT C4, INIT
C2834017|T037|S14.147A|ICD10CM|BROWN-SEQUARD SYNDROME AT C7 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|BROWN-SEQUARD SYNDROME AT C7, INIT
C2858886|T037|S72.463B|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL SUPRCNDL FX W INTRCNDL EXTN LOW END UNSP FEMR, 7THB
C2858887|T037|S72.463C|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL SUPRCNDL FX W INTRCNDL EXTN LOW END UNSP FEMR, 7THC
C2834045|T037|S14.154D|ICD10CM|OTHER INCOMPLETE LESION AT C4 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|OTH INCOMPLETE LESION AT C4, SUBS
C2875308|T046||ICD10CM|SEQUELAE OF GUILLAIN-BARRE SYNDROME
C2875309|T046|G65.1|ICD10CM|SEQUELAE OF OTHER INFLAMMATORY POLYNEUROPATHY|SEQUELAE OF OTHER INFLAMMATORY POLYNEUROPATHY
C2875310|T046||ICD10CM|SEQUELAE OF TOXIC POLYNEUROPATHY
C2890739|T037|T84.296A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTERNAL FIXATION DEVICE OF VERTEBRAE, INITIAL ENCOUNTER|MECH COMPL OF INTERNAL FIXATION DEVICE OF VERTEBRAE, INIT
C2832555|T037|S06.811S|ICD10CM|INJURY OF RIGHT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|INJ R INT CRTD, INTCR W LOC OF 30 MINUTES OR LESS, SEQUELA
C2832672|T037|S06.9X0A|ICD10CM|UNSPECIFIED INTRACRANIAL INJURY WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|UNSP INTRACRANIAL INJURY W/O LOSS OF CONSCIOUSNESS, INIT
C2887449|T047||ICD10CM|MILD INTERMITTENT ASTHMA, UNCOMPLICATED
C2887450|T047|J45.21|ICD10CM|MILD INTERMITTENT ASTHMA WITH (ACUTE) EXACERBATION|MILD INTERMITTENT ASTHMA WITH (ACUTE) EXACERBATION
C2887451|T047|J45.22|ICD10CM|MILD INTERMITTENT ASTHMA WITH STATUS ASTHMATICUS|MILD INTERMITTENT ASTHMA WITH STATUS ASTHMATICUS
C2977015|T047|I82.5Z1|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF RIGHT DISTAL LOWER EXTREMITY|CHR EMBLSM AND THOMBOS UNSP DEEP VEINS OF R DIST LOW EXTRM
C2977016|T047|I82.5Z2|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF LEFT DISTAL LOWER EXTREMITY|CHR EMBLSM AND THOMBOS UNSP DEEP VN OF LEFT DIST LOW EXTRM
C2977017|T047|I82.5Z3|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF DISTAL LOWER EXTREMITY, BILATERAL|CHR EMBLSM AND THOMBOS UNSP DEEP VEINS OF DIST LOW EXTRM, BI
C2977018|T047|I82.5Z9|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF UNSPECIFIED DISTAL LOWER EXTREMITY|CHR EMBLSM AND THOMBOS UNSP DEEP VN UNSP DISTAL LOW EXTRM
C2869820|T037|S98.141A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF ONE RIGHT LESSER TOE, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF ONE RIGHT LESSER TOE, INIT
C2882990|T047|I70.729|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, UNSPECIFIED EXTREMITY|ATHSCL TYPE OF BYPASS OF THE EXTRM W REST PAIN, UNSP EXTRM
C2882989|T047|I70.728|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, OTHER EXTREMITY|ATHSCL TYPE OF BYPASS OF THE EXTRM W REST PAIN, OTH EXTRM
C2882988|T047|I70.723|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, BILATERAL LEGS|ATHSCL TYPE OF BYPASS OF THE EXTRM W REST PAIN, BI LEGS
C2882987|T047|I70.722|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, LEFT LEG|ATHSCL TYPE OF BYPASS OF THE EXTRM W REST PAIN, LEFT LEG
C2882986|T047|I70.721|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, RIGHT LEG|ATHSCL TYPE OF BYPASS OF THE EXTRM W REST PAIN, RIGHT LEG
C2845936|T191|C72.41|ICD10CM|MALIGNANT NEOPLASM OF RIGHT ACOUSTIC NERVE|MALIGNANT NEOPLASM OF RIGHT ACOUSTIC NERVE
C2845935|T191|C72.40|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED ACOUSTIC NERVE|MALIGNANT NEOPLASM OF UNSPECIFIED ACOUSTIC NERVE
C2845937|T191|C72.42|ICD10CM|MALIGNANT NEOPLASM OF LEFT ACOUSTIC NERVE|MALIGNANT NEOPLASM OF LEFT ACOUSTIC NERVE
C2888909|T047|M00.841|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, RIGHT HAND|ARTHRITIS DUE TO OTHER BACTERIA, RIGHT HAND
C2888910|T047|M00.842|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, LEFT HAND|ARTHRITIS DUE TO OTHER BACTERIA, LEFT HAND
C2888911|T047|M00.849|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, UNSPECIFIED HAND|ARTHRITIS DUE TO OTHER BACTERIA, UNSPECIFIED HAND
C2834019|T037|S14.147S|ICD10CM|BROWN-SEQUARD SYNDROME AT C7 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|BROWN-SEQUARD SYNDROME AT C7, SEQUELA
C2893646|T047|M12.059|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], UNSPECIFIED HIP|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], UNSPECIFIED HIP
C2890513|T037|T84.052A|ICD10CM|PERIPROSTHETIC OSTEOLYSIS OF INTERNAL PROSTHETIC RIGHT KNEE JOINT, INITIAL ENCOUNTER|PERIPROSTH OSTEOLYSIS OF INTERNAL PROSTHETIC R KNEE JT, INIT
C4269452|T037|S02.611S|ICD10CM|FRACTURE OF CONDYLAR PROCESS OF RIGHT MANDIBLE, SEQUELA|FRACTURE OF CONDYLAR PROCESS OF RIGHT MANDIBLE, SEQUELA
C2882930|T047|I70.622|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, LEFT LEG|ATHSCL NONBIOL BYPASS OF THE EXTRM W REST PAIN, LEFT LEG
C2882931|T047|I70.623|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, BILATERAL LEGS|ATHSCL NONBIOL BYPASS OF THE EXTRM W REST PAIN, BI LEGS
C0260984|T067|E802.0|ICD9CM|UNSPECIFIED PORPHYRIA|RR ACC W DERAIL-EMPLOYEE
C2882929|T047|I70.621|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, RIGHT LEG|ATHSCL NONBIOL BYPASS OF THE EXTRM W REST PAIN, RIGHT LEG
C2874680|T048||ICD10CM|HALLUCINOGEN ABUSE WITH INTOXICATION, UNCOMPLICATED
C2874681|T048|F16.121|ICD10CM|HALLUCINOGEN ABUSE WITH INTOXICATION WITH DELIRIUM|HALLUCINOGEN ABUSE WITH INTOXICATION WITH DELIRIUM
C2874682|T048|F16.122|ICD10CM|HALLUCINOGEN ABUSE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE|HALLUCINOGEN ABUSE W INTOXICATION W PERCEPTUAL DISTURBANCE
C2832553|T037|S06.811A|ICD10CM|INJURY OF RIGHT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|INJ R INT CAROTID, INTCR W LOC OF 30 MINUTES OR LESS, INIT
C2886396|T037|T71.152S|ICD10CM|ASPHYXIATION DUE TO SMOTHERING IN FURNITURE, INTENTIONAL SELF-HARM, SEQUELA|ASPHYX DUE TO SMOTHERING IN FURNITURE, SELF-HARM, SEQUELA
C2882932|T047|I70.628|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, OTHER EXTREMITY|ATHSCL NONBIOL BYPASS OF THE EXTRM W REST PAIN, OTH EXTRM
C2882933|T047|I70.629|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, UNSPECIFIED EXTREMITY|ATHSCL NONBIOL BYPASS OF THE EXTRM W REST PAIN, UNSP EXTRM
C2874683|T048|F16.129|ICD10CM|HALLUCINOGEN ABUSE WITH INTOXICATION, UNSPECIFIED|HALLUCINOGEN ABUSE WITH INTOXICATION, UNSPECIFIED
C2901039|T046|M84.463A|ICD10CM|PATHOLOGICAL FRACTURE, RIGHT FIBULA, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, RIGHT FIBULA, INIT FOR FX
C2833399|T037|S12.330B|ICD10CM|UNSPECIFIED TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP TRAUM DISPL SPONDYLOLYSIS OF 4TH CERVCAL VERT, 7THB
C2833398|T037|S12.330A|ICD10CM|UNSPECIFIED TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP TRAUM DISPL SPONDYLOLYSIS OF FOURTH CERVCAL VERT, INIT
C2890666|T037|T84.192A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTERNAL FIXATION DEVICE OF BONE OF RIGHT FOREARM, INITIAL ENCOUNTER|MECH COMPL OF INT FIX OF BONE OF RIGHT FOREARM, INIT
C0153446|T191|C21.0|DMDICD10|MALIGNANT NEOPLASM OF ANUS, UNSPECIFIED|BOESARTIGE NEUBILDUNG: ANUS, NICHT NAEHER BEZEICHNET
C0864874|T191||ICD10CM|MALIGNANT NEOPLASM OF ANAL CANAL
C0345886|T191|C21.2|DMDICD10|MALIGNANT NEOPLASM OF CLOACOGENIC ZONE|BOESARTIGE NEUBILDUNG: KLOAKENREGION
C2837937|T191|C21.8|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF RECTUM, ANUS AND ANAL CANAL|PRIMARY MALIGNANT NEOPLASM OF TWO OR MORE CONTIGUOUS SITES OF RECTUM, ANUS AND ANAL CANAL
C2883785|T037|T50.992A|ICD10CM|POISONING BY OTHER DRUGS, MEDICAMENTS AND BIOLOGICAL SUBSTANCES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH DRUG/MEDS/BIOL SUBST, SELF-HARM, INIT
C2832475|T037|S06.5X1S|ICD10CM|TRAUMATIC SUBDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|TRAUM SUBDR HEM W LOC OF 30 MINUTES OR LESS, SEQUELA
C2832230|T037|S06.342S|ICD10CM|TRAUMATIC HEMORRHAGE OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|TRAUM HEMOR RIGHT CEREBRUM W LOC OF 31-59 MIN, SEQUELA
C4509334|T047|L97.918|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF RIGHT LOWER LEG WITH OTHER SPECIFIED SEVERITY|NON-PRS CHRONIC ULC UNSP PRT OF R LOW LEG WITH OTH SEVERITY
C2888765|T047|L97.919|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF RIGHT LOWER LEG WITH UNSPECIFIED SEVERITY|NON-PRS CHRONIC ULC UNSP PRT OF R LOW LEG W UNSP SEVERITY
C2891001|T037|T85.199A|ICD10CM|OTHER MECHANICAL COMPLICATION OF OTHER IMPLANTED ELECTRONIC STIMULATOR OF NERVOUS SYSTEM, INITIAL ENCOUNTER|MECH COMPL OF IMPLNT ELECTRNC STIMULTR OF NERVOUS SYS, INIT
C4270485|T046|T85.122A|ICD10CM|DISPLACEMENT OF IMPLANTED ELECTRONIC NEUROSTIMULATOR OF SPINAL CORD ELECTRODE (LEAD), INITIAL ENCOUNTER|DISPLACEMENT OF IMPLNT ELEC NSTIM OF SPINAL CORD LEAD, INIT
C2832473|T037|S06.5X1A|ICD10CM|TRAUMATIC SUBDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|TRAUM SUBDR HEM W LOC OF 30 MINUTES OR LESS, INIT
C2832228|T037|S06.342A|ICD10CM|TRAUMATIC HEMORRHAGE OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|TRAUM HEMOR RIGHT CEREBRUM W LOC OF 31-59 MIN, INIT
C2888761|T047|L97.911|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF RIGHT LOWER LEG LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHR ULC UNSP PRT OF R LOW LEG LIMITED TO BRKDWN SKIN
C2888762|T047|L97.912|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF RIGHT LOWER LEG WITH FAT LAYER EXPOSED|NON-PRS CHR ULC UNSP PRT OF R LOW LEG W FAT LAYER EXPOSED
C2888763|T047|L97.913|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF RIGHT LOWER LEG WITH NECROSIS OF MUSCLE|NON-PRS CHRONIC ULC UNSP PRT OF R LOW LEG W NECROS MUSCLE
C2888764|T047|L97.914|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF RIGHT LOWER LEG WITH NECROSIS OF BONE|NON-PRS CHRONIC ULC UNSP PRT OF R LOW LEG W NECROSIS OF BONE
C4509332|T047|L97.915|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF RIGHT LOWER LEG WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC UNSP PRT R LW LEG W MSL INVL W/O EVD OF NECR
C4509333|T047|L97.916|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF RIGHT LOWER LEG WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC UNSP PRT R LW LEG W BNE INVL W/O EVD OF NECR
C2900490|T047|B01.12|ICD10CM|VARICELLA MYELITIS|VARICELLA MYELITIS
C2833643|T037|S12.691A|ICD10CM|OTHER NONDISPLACED FRACTURE OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH NONDISP FX OF SEVENTH CERVICAL VERTEBRA, INIT
C2833644|T037|S12.691B|ICD10CM|OTHER NONDISPLACED FRACTURE OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH NONDISP FX OF SEVENTH CERVICAL VERTEBRA, INIT FOR OPN FX
C0042909|T046|H43.10|ICD10CM|VITREOUS HEMORRHAGE, UNSPECIFIED EYE|VITREOUS HEMORRHAGE, UNSPECIFIED EYE
C2833146|T037|S12.001B|ICD10CM|UNSPECIFIED NONDISPLACED FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP NONDISP FX OF FIRST CERVICAL VERTEBRA, INIT FOR OPN FX
C2832111|T037|S06.314A|ICD10CM|CONTUSION AND LACERATION OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|CONTUS/LAC RIGHT CEREBRUM W LOC OF 6 HOURS TO 24 HOURS, INIT
C4268162|T047|E13.3539|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, UNSPECIFIED EYE|OTH DIAB WITH PROLIF DIAB RTNOP WITH TRCTN DTCH N-MCLA, UNSP
C2888787|T047|L98.491|ICD10CM|NON-PRESSURE CHRONIC ULCER OF SKIN OF OTHER SITES LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHRONIC ULCER SKIN/ SITES LIMITED TO BRKDWN SKIN
C2888788|T047|L98.492|ICD10CM|NON-PRESSURE CHRONIC ULCER OF SKIN OF OTHER SITES WITH FAT LAYER EXPOSED|NON-PRS CHRONIC ULCER OF SKIN OF SITES W FAT LAYER EXPOSED
C2888789|T047|L98.493|ICD10CM|NON-PRESSURE CHRONIC ULCER OF SKIN OF OTHER SITES WITH NECROSIS OF MUSCLE|NON-PRS CHRONIC ULCER OF SKIN OF SITES W NECROSIS OF MUSCLE
C2888790|T047|L98.494|ICD10CM|NON-PRESSURE CHRONIC ULCER OF SKIN OF OTHER SITES WITH NECROSIS OF BONE|NON-PRS CHRONIC ULCER OF SKIN OF SITES W NECROSIS OF BONE
C4509344|T047|L98.495|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER SITES WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULCER OF SITES WITH MUSCLE INVL W/O EVD OF NECR
C4509345|T047|L98.496|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER SITES WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULCER OF SITES WITH BONE INVL W/O EVD OF NECR
C4509346|T047|L98.498|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER SITES WITH OTHER SPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF OTHER SITES WITH OTH SEVERITY
C2888791|T047|L98.499|ICD10CM|NON-PRESSURE CHRONIC ULCER OF SKIN OF OTHER SITES WITH UNSPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF SKIN OF SITES W UNSP SEVERITY
C2901929|T047|M86.662|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, LEFT TIBIA AND FIBULA|OTHER CHRONIC OSTEOMYELITIS, LEFT TIBIA AND FIBULA
C2901928|T047|M86.661|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, RIGHT TIBIA AND FIBULA|OTHER CHRONIC OSTEOMYELITIS, RIGHT TIBIA AND FIBULA
C2835859|T037|S24.159S|ICD10CM|OTHER INCOMPLETE LESION AT UNSPECIFIED LEVEL OF THORACIC SPINAL CORD, SEQUELA|OTH INCMPL LESION AT UNSP LEVEL OF THOR SPINAL CORD, SEQUELA
C2873990|T047|E09.49|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH NEUROLOGICAL COMPLICATIONS WITH OTHER DIABETIC NEUROLOGICAL COMPLICATION|DRUG/CHEM DIABETES W NEURO COMP W OTH DIABETIC NEURO COMP
C2842092|T191|C50.212|ICD10CM|MALIGNANT NEOPLASM OF UPPER-INNER QUADRANT OF LEFT FEMALE BREAST|MALIG NEOPLASM OF UPPER-INNER QUADRANT OF LEFT FEMALE BREAST
C2842091|T191|C50.211|ICD10CM|MALIGNANT NEOPLASM OF UPPER-INNER QUADRANT OF RIGHT FEMALE BREAST|MALIG NEOPLM OF UPPER-INNER QUADRANT OF RIGHT FEMALE BREAST
C2873989|T047|E09.44|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH NEUROLOGICAL COMPLICATIONS WITH DIABETIC AMYOTROPHY|DRUG/CHEM DIABETES W NEUROLOGICAL COMP W DIABETIC AMYOTROPHY
C4267980|T047|E09.3513|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|DRUG/CHEM DIAB WITH PROLIF DIAB RTNOP WITH MACULAR EDEMA, BI
C2842152|T191|C57.11|ICD10CM|MALIGNANT NEOPLASM OF RIGHT BROAD LIGAMENT|MALIGNANT NEOPLASM OF RIGHT BROAD LIGAMENT
C2842151|T191|C57.10|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED BROAD LIGAMENT|MALIGNANT NEOPLASM OF UNSPECIFIED BROAD LIGAMENT
C2842093|T191|C50.219|ICD10CM|MALIGNANT NEOPLASM OF UPPER-INNER QUADRANT OF UNSPECIFIED FEMALE BREAST|MALIG NEOPLASM OF UPPER-INNER QUADRANT OF UNSP FEMALE BREAST
C2842153|T191|C57.12|ICD10CM|MALIGNANT NEOPLASM OF LEFT BROAD LIGAMENT|MALIGNANT NEOPLASM OF LEFT BROAD LIGAMENT
C2876868|T037|T37.3X2A|ICD10CM|POISONING BY OTHER ANTIPROTOZOAL DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH ANTIPROTOZOAL DRUGS, SELF-HARM, INIT
C2885767|T037|T63.612S|ICD10CM|TOXIC EFFECT OF CONTACT WITH PORTUGESE MAN-O-WAR, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CNTCT W PORTUGESE MAN-O-WAR, SLF-HRM, SQLA
C0836987|T047||ICD10CM|TYPE 1 DIABETES MELLITUS WITH KETOACIDOSIS WITHOUT COMA
C0836988|T047||ICD10CM|TYPE 1 DIABETES MELLITUS WITH KETOACIDOSIS WITH COMA
C2882707|T047|I70.228|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES WITH REST PAIN, OTHER EXTREMITY|ATHSCL NATIVE ARTERIES OF EXTRM W REST PAIN, OTH EXTREMITY
C0432420|T047|Q91.2|DMDICD10|TRISOMY 18, TRANSLOCATION|TRISOMIE 18, TRANSLOKATION
C0432426|T049|Q91.5|DMDICD10|TRISOMY 13, MOSAICISM (MITOTIC NONDISJUNCTION)|TRISOMIE 13, MOSAIK (MITOTISCHE NON-DISJUNCTION)
C2910355|T047||ICD10CM|TRISOMY 13, NONMOSAICISM (MEIOTIC NONDISJUNCTION)
C0152095|T047|Q91.7|DMDICD10|TRISOMY 13, UNSPECIFIED|PATAU-SYNDROM, NICHT NAEHER BEZEICHNET
C0432424|T047|Q91.6|DMDICD10|TRISOMY 13, TRANSLOCATION|TRISOMIE 13, TRANSLOKATION
C2919144|T191|C19|ICD10CM|MALIGNANT NEOPLASM OF RECTOSIGMOID JUNCTION|MALIGNANT NEOPLASM OF COLON WITH RECTUM
C0153400|T191|C12|DMDICD10|MALIGNANT NEOPLASM OF PYRIFORM SINUS|BOESARTIGE NEUBILDUNG DES RECESSUS PIRIFORMIS
C4270276|T046|T83.193A|ICD10CM|OTHER MECHANICAL COMPLICATION OF OTHER URINARY STENT, INITIAL ENCOUNTER|MECH COMPL OF OTHER URINARY STENT, INITIAL ENCOUNTER
C2860149|T037|S79.112A|ICD10CM|SALTER-HARRIS TYPE I PHYSEAL FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SLTR-HARIS TYPE I PHYSEAL FX LOWER END OF LEFT FEMUR, INIT
C2858303|T037|S72.402A|ICD10CM|UNSPECIFIED FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF LOWER END OF LEFT FEMUR, INIT FOR CLOS FX
C2858305|T037|S72.402C|ICD10CM|UNSPECIFIED FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP FX LOWER END OF LEFT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2858304|T037|S72.402B|ICD10CM|UNSPECIFIED FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP FX LOWER END OF LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C0153290|T047|B67.1|DMDICD10|ECHINOCOCCUS GRANULOSUS INFECTION OF LUNG|ECHINOCOCCUS-GRANULOSUS-INFEKTION [ZYSTISCHE ECHINOKOKKOSE] DER LUNGE
C2873779|T047|D61.89|ICD10CM|OTHER SPECIFIED APLASTIC ANEMIAS AND OTHER BONE MARROW FAILURE SYNDROMES|OTH APLASTIC ANEMIAS AND OTHER BONE MARROW FAILURE SYNDROMES
C0302112|T047|D61.82|ICD10CM|MYELOPHTHISIS|MYELOPHTHISIS
C2883912|T037|T50.B92A|ICD10CM|POISONING BY OTHER VIRAL VACCINES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH VIRAL VACCINES, INTENTIONAL SELF-HARM, INIT
C2837783|T037|S32.17XB|ICD10CM|TYPE 4 FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE 4 FRACTURE OF SACRUM, INIT ENCNTR FOR OPEN FRACTURE
C2837782|T037|S32.17XA|ICD10CM|TYPE 4 FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE 4 FRACTURE OF SACRUM, INIT ENCNTR FOR CLOSED FRACTURE
C2960068|T191|C49.A4|ICD10CM|GASTROINTESTINAL STROMAL TUMOR OF LARGE INTESTINE|GASTROINTESTINAL STROMAL TUMOR OF LARGE INTESTINE
C4267835|T191|C49.A5|ICD10CM|GASTROINTESTINAL STROMAL TUMOR OF RECTUM|GASTROINTESTINAL STROMAL TUMOR OF RECTUM
C2883914|T037|T50.B92S|ICD10CM|POISONING BY OTHER VIRAL VACCINES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH VIRAL VACCINES, SELF-HARM, SEQUELA
C4267834|T191|C49.A0|ICD10CM|GASTROINTESTINAL STROMAL TUMOR, UNSPECIFIED SITE|GASTROINTESTINAL STROMAL TUMOR, UNSPECIFIED SITE
C2959942|T191|C49.A1|ICD10CM|GASTROINTESTINAL STROMAL TUMOR OF ESOPHAGUS|GASTROINTESTINAL STROMAL TUMOR OF ESOPHAGUS
C1333768|T191|C49.A2|ICD10CM|GASTROINTESTINAL STROMAL TUMOR OF STOMACH|GASTROINTESTINAL STROMAL TUMOR OF STOMACH
C1335996|T191|C49.A3|ICD10CM|GASTROINTESTINAL STROMAL TUMOR OF SMALL INTESTINE|GASTROINTESTINAL STROMAL TUMOR OF SMALL INTESTINE
C4267836|T191|C49.A9|ICD10CM|GASTROINTESTINAL STROMAL TUMOR OF OTHER SITES|GASTROINTESTINAL STROMAL TUMOR OF OTHER SITES
C0014065|T019|Q01.9|DMDICD10|ENCEPHALOCELE, UNSPECIFIED|ENZEPHALOZELE, NICHT NAEHER BEZEICHNET
C1142536|T047||ICD10CM|PNEUMONIA DUE TO METHICILLIN RESISTANT STAPHYLOCOCCUS AUREUS
C2349530|T047||ICD10CM|PNEUMONIA DUE TO METHICILLIN SUSCEPTIBLE STAPHYLOCOCCUS AUREUS
C2889980|T037|T82.41XS|ICD10CM|BREAKDOWN (MECHANICAL) OF VASCULAR DIALYSIS CATHETER, SEQUELA|BREAKDOWN OF VASCULAR DIALYSIS CATHETER, SEQUELA
C2860097|T037|S79.091A|ICD10CM|OTHER PHYSEAL FRACTURE OF UPPER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH PHYSEAL FRACTURE OF UPPER END OF RIGHT FEMUR, INIT
C2889535|T047|M08.041|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, RIGHT HAND|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, RIGHT HAND
C2889536|T047|M08.042|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, LEFT HAND|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, LEFT HAND
C2889979|T037|T82.41XD|ICD10CM|BREAKDOWN (MECHANICAL) OF VASCULAR DIALYSIS CATHETER, SUBSEQUENT ENCOUNTER|BREAKDOWN (MECHANICAL) OF VASCULAR DIALYSIS CATHETER, SUBS
C2889537|T047|M08.04|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED HAND|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, HAND
C2889978|T037|T82.41XA|ICD10CM|BREAKDOWN (MECHANICAL) OF VASCULAR DIALYSIS CATHETER, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF VASCULAR DIALYSIS CATHETER, INIT
C2890546|T037|T84.068A|ICD10CM|WEAR OF ARTICULAR BEARING SURFACE OF OTHER INTERNAL PROSTHETIC JOINT, INITIAL ENCOUNTER|WEAR OF ARTIC BEARING SURFACE OF INTERNAL PROSTH JOINT, INIT
C2858096|T037|S72.355A|ICD10CM|NONDISPLACED COMMINUTED FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP COMMINUTED FRACTURE OF SHAFT OF LEFT FEMUR, INIT
C2858097|T037|S72.355B|ICD10CM|NONDISPLACED COMMINUTED FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP COMMNT FX SHAFT OF L FEMUR, INIT FOR OPN FX TYPE I/2
C2858098|T037|S72.355C|ICD10CM|NONDISPLACED COMMINUTED FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP COMMNT FX SHAFT OF L FEMR, 7THC
C2843292|T037|S48.029S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT UNSPECIFIED SHOULDER JOINT, SEQUELA|PARTIAL TRAUMATIC AMPUTATION AT UNSP SHOULDER JOINT, SEQUELA
C2856023|T037|S68.615S|ICD10CM|COMPLETE TRAUMATIC TRANSPHALANGEAL AMPUTATION OF LEFT RING FINGER, SEQUELA|COMPLETE TRAUMATIC TRNSPHAL AMP OF L RNG FNGR, SEQUELA
C0375735|T067|E880.1|ICD9CM|ALPHA-1-ANTITRYPSIN DEFICIENCY|FALL ON SIDEWALK CURB
C2889113|T047|M05.022|ICD10CM|FELTY'S SYNDROME, LEFT ELBOW|FELTY'S SYNDROME, LEFT ELBOW
C4270573|T046|T85.731A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO IMPLANTED ELECTRONIC NEUROSTIMULATOR OF BRAIN, ELECTRODE (LEAD), INITIAL ENCOUNTER|I/I REACT D/T IMPLNT ELEC NSTIM OF BRAIN, LEAD, INIT
C3469320|T047|M05.029|ICD10CM|FELTY'S SYNDROME, UNSPECIFIED ELBOW|FELTY'S SYNDROME, UNSPECIFIED ELBOW
C2886017|T037|T65.212S|ICD10CM|TOXIC EFFECT OF CHEWING TOBACCO, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CHEWING TOBACCO, SELF-HARM, SEQUELA
C2845907|T191|C69.22|ICD10CM|MALIGNANT NEOPLASM OF LEFT RETINA|MALIGNANT NEOPLASM OF LEFT RETINA
C2837948|T191|C34.01|ICD10CM|MALIGNANT NEOPLASM OF RIGHT MAIN BRONCHUS|MALIGNANT NEOPLASM OF RIGHT MAIN BRONCHUS
C2845905|T191|C69.20|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED RETINA|MALIGNANT NEOPLASM OF UNSPECIFIED RETINA
C2888953|T047|M01.X69|ICD10CM|DIRECT INFECTION OF UNSPECIFIED KNEE IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIRECT INFCT OF UNSP KNEE IN INFEC/PARASTC DIS CLASSD ELSWHR
C2882373|T047|I63.332|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF LEFT POSTERIOR CEREBRAL ARTERY|CEREBRAL INFRC DUE TO THOMBOS OF LEFT POST CEREBRAL ARTERY
C2886015|T037|T65.212A|ICD10CM|TOXIC EFFECT OF CHEWING TOBACCO, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CHEWING TOBACCO, INTENTIONAL SELF-HARM, INIT
C2888951|T047|M01.X61|ICD10CM|DIRECT INFECTION OF RIGHT KNEE IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIRECT INFCT OF R KNEE IN INFEC/PARASTC DIS CLASSD ELSWHR
C2888952|T047|M01.X62|ICD10CM|DIRECT INFECTION OF LEFT KNEE IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIRECT INFCT OF L KNEE IN INFEC/PARASTC DIS CLASSD ELSWHR
C2832571|T037|S06.815S|ICD10CM|INJURY OF RIGHT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, SEQUELA|INJ R INT CRTD, INTCR W LOC >24 HR W RET CONSC LEV, SEQUELA
C2832569|T037|S06.815A|ICD10CM|INJURY OF RIGHT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, INITIAL ENCOUNTER|INJ R INT CAROTID, INTCR W LOC >24 HR W RET CONSC LEV, INIT
C2856040|T037|S68.619S|ICD10CM|COMPLETE TRAUMATIC TRANSPHALANGEAL AMPUTATION OF UNSPECIFIED FINGER, SEQUELA|COMPLETE TRAUMATIC TRNSPHAL AMP OF UNSP FINGER, SEQUELA
C0153425|T191|C17.9|DMDICD10|MALIGNANT NEOPLASM OF SMALL INTESTINE, UNSPECIFIED|BOESARTIGE NEUBILDUNG: DUENNDARM, NICHT NAEHER BEZEICHNET
C0349050|T191|C17.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF SMALL INTESTINE|BOESARTIGE NEUBILDUNG: DUENNDARM, MEHRERE TEILBEREICHE UEBERLAPPEND
C0153427|T191|C17.1|DMDICD10|MALIGNANT NEOPLASM OF JEJUNUM|BOESARTIGE NEUBILDUNG: JEJUNUM
C0153426|T191|C17.0|DMDICD10|MALIGNANT NEOPLASM OF DUODENUM|BOESARTIGE NEUBILDUNG: DUODENUM
C2979886|T191|C17.3|ICD10CM|MECKEL'S DIVERTICULUM, MALIGNANT|MECKEL'S DIVERTICULUM, MALIGNANT
C0153428|T191|C17.2|DMDICD10|MALIGNANT NEOPLASM OF ILEUM|BOESARTIGE NEUBILDUNG: ILEUM
C2890422|T037|T84.019A|ICD10CM|BROKEN INTERNAL JOINT PROSTHESIS, UNSPECIFIED SITE, INITIAL ENCOUNTER|BROKEN INTERNAL JOINT PROSTHESIS, UNSP SITE, INIT ENCNTR
C2901314|T046|M84.571A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, RIGHT ANKLE, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, RIGHT ANKLE, INIT
C2902900|T047|N05.5|ICD10CM|UNSPECIFIED NEPHRITIC SYNDROME WITH DIFFUSE MESANGIOCAPILLARY GLOMERULONEPHRITIS|UNSPECIFIED NEPHRITIC SYNDROME WITH MEMBRANOPROLIFERATIVE GLOMERULONEPHRITIS, TYPES 1 AND 3, OR NOS
C0477723|T047|N05.4|DMDICD10|UNSPECIFIED NEPHRITIC SYNDROME WITH DIFFUSE ENDOCAPILLARY PROLIFERATIVE GLOMERULONEPHRITIS|NICHT NAEHER BEZEICHNETES NEPHRITISCHES SYNDROM: DIFFUSE ENDOKAPILLAER-PROLIFERATIVE GLOMERULONEPHRITIS
C2902902|T047|N05.7|ICD10CM|UNSPECIFIED NEPHRITIC SYNDROME WITH DIFFUSE CRESCENTIC GLOMERULONEPHRITIS|UNSPECIFIED NEPHRITIC SYNDROME WITH EXTRACAPILLARY GLOMERULONEPHRITIS
C0477377|T047|G46.8|DMDICD10|OTHER VASCULAR SYNDROMES OF BRAIN IN CEREBROVASCULAR DISEASES|SONSTIGE SYNDROME DER HIRNGEFAESSE BEI ZEREBROVASKULAEREN KRANKHEITEN
C2875088|T047|G40.119|ICD10CM|LOCALIZATION-RELATED (FOCAL) (PARTIAL) SYMPTOMATIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SIMPLE PARTIAL SEIZURES, INTRACTABLE, WITHOUT STATUS EPILEPTICUS|LOCAL-REL SYMPTC EPI W SIMPLE PART SEIZ, NTRCT, W/O STAT EPI
C2902896|T047|N05.0|ICD10CM|UNSPECIFIED NEPHRITIC SYNDROME WITH MINOR GLOMERULAR ABNORMALITY|UNSPECIFIED NEPHRITIC SYNDROME WITH MINIMAL CHANGE LESION
C0477722|T047|N05.3|DMDICD10|UNSPECIFIED NEPHRITIC SYNDROME WITH DIFFUSE MESANGIAL PROLIFERATIVE GLOMERULONEPHRITIS|NICHT NAEHER BEZEICHNETES NEPHRITISCHES SYNDROM: DIFFUSE MESANGIOPROLIFERATIVE GLOMERULONEPHRITIS
C0495032|T047|N05.2|DMDICD10|UNSPECIFIED NEPHRITIC SYNDROME WITH DIFFUSE MEMBRANOUS GLOMERULONEPHRITIS|NICHT NAEHER BEZEICHNETES NEPHRITISCHES SYNDROM: DIFFUSE MEMBRANOESE GLOMERULONEPHRITIS
C0455717|T047||ICD10CM|BRAIN STEM STROKE SYNDROME
C0451681|T047|G46.2|DMDICD10|POSTERIOR CEREBRAL ARTERY SYNDROME|ARTERIA-CEREBRI-POSTERIOR-SYNDROM
C0451680|T047|G46.1|DMDICD10|ANTERIOR CEREBRAL ARTERY SYNDROME|ARTERIA-CEREBRI-ANTERIOR-SYNDROM
C0238281|T047|G46.0|DMDICD10|MIDDLE CEREBRAL ARTERY SYNDROME|ARTERIA-CEREBRI-MEDIA-SYNDROM
C2875087|T047|G40.111|ICD10CM|LOCALIZATION-RELATED (FOCAL) (PARTIAL) SYMPTOMATIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SIMPLE PARTIAL SEIZURES, INTRACTABLE, WITH STATUS EPILEPTICUS|LOCAL-REL SYMPTC EPI W SIMPLE PART SEIZ, NTRCT, W STAT EPI
C0393958|T047|G46.6|DMDICD10|PURE SENSORY LACUNAR SYNDROME|REIN SENSORISCHES LAKUNAERES SYNDROM
C0393957|T047|G46.5|DMDICD10|PURE MOTOR LACUNAR SYNDROME|REIN MOTORISCHES LAKUNAERES SYNDROM
C0451672|T047|G46.4|DMDICD10|CEREBELLAR STROKE SYNDROME|KLEINHIRNSYNDROM
C2835227|T037|S22.020B|ICD10CM|WEDGE COMPRESSION FRACTURE OF SECOND THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|WEDGE COMPRSN FX SECOND THOR VERTEBRA, INIT FOR OPN FX
C2835226|T037|S22.020A|ICD10CM|WEDGE COMPRESSION FRACTURE OF SECOND THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|WEDGE COMPRESSION FRACTURE OF SECOND THORACIC VERTEBRA, INIT
C0152491|T047|A02.24|ICD10CM|SALMONELLA OSTEOMYELITIS|SALMONELLA OSTEOMYELITIS
C2905794|T037|X82.1XXA|ICD10CM|INTENTIONAL COLLISION OF MOTOR VEHICLE WITH TRAIN, INITIAL ENCOUNTER|INTENTIONAL COLLISION OF MOTOR VEHICLE W TRAIN, INIT ENCNTR
C0152489|T047|A02.22|ICD10CM|SALMONELLA PNEUMONIA|SALMONELLA PNEUMONIA
C0152490|T047|A02.23|ICD10CM|SALMONELLA ARTHRITIS|SALMONELLA ARTHRITIS
C2857205|T037|S72.114A|ICD10CM|NONDISPLACED FRACTURE OF GREATER TROCHANTER OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF GREATER TROCHANTER OF RIGHT FEMUR, INIT
C0043046|T047||ICD10CM|CACHEXIA
C2905796|T037|X82.1XXS|ICD10CM|INTENTIONAL COLLISION OF MOTOR VEHICLE WITH TRAIN, SEQUELA|INTENTIONAL COLLISION OF MOTOR VEHICLE WITH TRAIN, SEQUELA
C2832146|T037|S06.322S|ICD10CM|CONTUSION AND LACERATION OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|CONTUS/LAC LEFT CEREBRUM W LOC OF 31-59 MIN, SEQUELA
C4267851|T191|C81.29|ICD10CM|MIXED CELLULARITY HODGKIN LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES|MIXED CELLULAR HODGKIN LYMPH, EXTRNOD AND SOLID ORGAN SITES
C4267850|T191|C81.28|ICD10CM|MIXED CELLULARITY HODGKIN LYMPHOMA, LYMPH NODES OF MULTIPLE SITES|MIXED CELLULARITY HODGKIN LYMPHOMA, LYMPH NODES MULT SITE
C2857206|T037|S72.114B|ICD10CM|NONDISPLACED FRACTURE OF GREATER TROCHANTER OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF GREATER TROCHANTER OF R FEMR, 7THB
C2896575|T046|M80.051A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, RIGHT FEMUR, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, RIGHT FEMUR, INIT
C2887484|T047|J80|ICD10CM|ACUTE RESPIRATORY DISTRESS SYNDROME|ACUTE RESPIRATORY DISTRESS SYNDROME IN ADULT OR CHILD
C0153768|T191|C81.21|ICD10CM|MIXED CELLULARITY HODGKIN LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK|MIXED CELLULAR HODGKIN LYMPH, NODES OF HEAD, FACE, AND NECK
C4267845|T191|C81.20|ICD10CM|MIXED CELLULARITY HODGKIN LYMPHOMA, UNSPECIFIED SITE|MIXED CELLULARITY HODGKIN LYMPHOMA, UNSPECIFIED SITE
C4267847|T191|C81.23|ICD10CM|MIXED CELLULARITY HODGKIN LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES|MIXED CELLULARITY HODGKIN LYMPHOMA, INTRA-ABD LYMPH NODES
C4267846|T191|C81.22|ICD10CM|MIXED CELLULARITY HODGKIN LYMPHOMA, INTRATHORACIC LYMPH NODES|MIXED CELLULARITY HODGKIN LYMPHOMA, INTRATHORAC LYMPH NODES
C4267848|T191|C81.25|ICD10CM|MIXED CELLULARITY HODGKIN LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|MIXED CELLULAR HDGKN LYMPH, NODES OF ING RGN AND LOWER LIMB
C0153771|T191|C81.24|ICD10CM|MIXED CELLULARITY HODGKIN LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB|MIXED CELLULAR HODGKIN LYMPH, NODES OF AXILLA AND UPPER LIMB
C0153774|T191||ICD10CM|MIXED CELLULARITY HODGKIN LYMPHOMA, SPLEEN
C2882881|T047|I70.533|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF ANKLE|ATHSCL NONAUT BIO BYPASS OF THE RIGHT LEG W ULCER OF ANKLE
C2888993|T047|M02.111|ICD10CM|POSTDYSENTERIC ARTHROPATHY, RIGHT SHOULDER|POSTDYSENTERIC ARTHROPATHY, RIGHT SHOULDER
C2888994|T047|M02.112|ICD10CM|POSTDYSENTERIC ARTHROPATHY, LEFT SHOULDER|POSTDYSENTERIC ARTHROPATHY, LEFT SHOULDER
C2838243|T037|S32.464A|ICD10CM|NONDISPLACED ASSOCIATED TRANSVERSE-POSTERIOR FRACTURE OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP ASSOCIATED TRANSV/POST FX RIGHT ACETABULUM, INIT
C2838244|T037|S32.464B|ICD10CM|NONDISPLACED ASSOCIATED TRANSVERSE-POSTERIOR FRACTURE OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP ASSOC TRANSV/POST FX RIGHT ACETAB, INIT FOR OPN FX
C2888995|T047|M02.119|ICD10CM|POSTDYSENTERIC ARTHROPATHY, UNSPECIFIED SHOULDER|POSTDYSENTERIC ARTHROPATHY, UNSPECIFIED SHOULDER
C2882879|T047|I70.531|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF THIGH|ATHSCL NONAUT BIO BYPASS OF THE RIGHT LEG W ULCER OF THIGH
C2891268|T037|T86.09|ICD10CM|OTHER COMPLICATIONS OF BONE MARROW TRANSPLANT|OTHER COMPLICATIONS OF BONE MARROW TRANSPLANT
C2859198|T037|S73.024A|ICD10CM|OBTURATOR DISLOCATION OF RIGHT HIP, INITIAL ENCOUNTER|OBTURATOR DISLOCATION OF RIGHT HIP, INITIAL ENCOUNTER
C2885697|T037|T63.462S|ICD10CM|TOXIC EFFECT OF VENOM OF WASPS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF WASPS, SELF-HARM, SEQUELA
C2891267|T046||ICD10CM|BONE MARROW TRANSPLANT INFECTION
C0340991|T046|T86.02|ICD10CM|BONE MARROW TRANSPLANT FAILURE|BONE MARROW TRANSPLANT FAILURE
C0340990|T046|T86.01|ICD10CM|BONE MARROW TRANSPLANT REJECTION|BONE MARROW TRANSPLANT REJECTION
C2891266|T037|T86.00|ICD10CM|UNSPECIFIED COMPLICATION OF BONE MARROW TRANSPLANT|UNSPECIFIED COMPLICATION OF BONE MARROW TRANSPLANT
C2874801|T048|F19.16|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE ABUSE WITH PSYCHOACTIVE SUBSTANCE-INDUCED PERSISTING AMNESTIC DISORDER|OTH PSYCHOACTV SUBSTANCE ABUSE W PERSIST AMNESTIC DISORDER
C4268286|T048|F19.17|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE ABUSE WITH PSYCHOACTIVE SUBSTANCE-INDUCED PERSISTING DEMENTIA|OTHER (OR UNKNOWN) SUBSTANCE USE DISORDER, MILD, WITH OTHER (OR UNKNOWN) SUBSTANCE-INDUCED MAJOR NEUROCOGNITIVE DISORDER
C4268285|T048|F19.14|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE ABUSE WITH PSYCHOACTIVE SUBSTANCE-INDUCED MOOD DISORDER|OTHER (OR UNKNOWN) SUBSTANCE USE DISORDER, MILD, WITH OTHER (OR UNKNOWN) SUBSTANCE-INDUCED DEPRESSIVE DISORDER
C2885695|T037|T63.462A|ICD10CM|TOXIC EFFECT OF VENOM OF WASPS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF WASPS, INTENTIONAL SELF-HARM, INIT
C2884931|T037|T59.6X2S|ICD10CM|TOXIC EFFECT OF HYDROGEN SULFIDE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF HYDROGEN SULFIDE, SELF-HARM, SEQUELA
C2874807|T048|F19.19|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE ABUSE WITH UNSPECIFIED PSYCHOACTIVE SUBSTANCE-INDUCED DISORDER|OTH PSYCHOACTIVE SUBSTANCE ABUSE W UNSP DISORDER
C4509596|T047|E85.4|ICD10CM|ORGAN-LIMITED AMYLOIDOSIS|TRANSTHYRETIN-RELATED (ATTR) FAMILIAL AMYLOID CARDIOMYOPATHY
C2874525|T048|F13.19|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE WITH UNSPECIFIED SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED DISORDER|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE W UNSP DISORDER
C2869875|T037|S98.321D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT MIDFOOT, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF RIGHT MIDFOOT, SUBS ENCNTR
C1719313|T047||ICD10CM|NON-NEUROPATHIC HEREDOFAMILIAL AMYLOIDOSIS
C4509022|T047|E85.1|ICD10CM|NEUROPATHIC HEREDOFAMILIAL AMYLOIDOSIS|TRANSTHYRETIN-RELATED (ATTR) FAMILIAL AMYLOID POLYNEUROPATHY
C0348506|T047|E85.2|DMDICD10|HEREDOFAMILIAL AMYLOIDOSIS, UNSPECIFIED|HEREDOFAMILIAERE AMYLOIDOSE, NICHT NAEHER BEZEICHNET
C3536716|T047|E85.3|DMDICD10|SECONDARY SYSTEMIC AMYLOIDOSIS|SEKUNDAERE SYSTEMISCHE AMYLOIDOSE
C2874478|T048|F12.151|ICD10CM|CANNABIS ABUSE WITH PSYCHOTIC DISORDER WITH HALLUCINATIONS|CANNABIS ABUSE WITH PSYCHOTIC DISORDER WITH HALLUCINATIONS
C2874477|T048|F12.150|ICD10CM|CANNABIS ABUSE WITH PSYCHOTIC DISORDER WITH DELUSIONS|CANNABIS ABUSE WITH PSYCHOTIC DISORDER WITH DELUSIONS
C2838172|T037|S32.446B|ICD10CM|NONDISPLACED FRACTURE OF POSTERIOR COLUMN [ILIOISCHIAL] OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP FX OF POST COLUMN OF UNSP ACETAB, INIT FOR OPN FX
C4268221|T048|F13.14|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED MOOD DISORDER|SEDATIVE, HYPNOTIC, OR ANXIOLYTIC USE DISORDER, MILD, WITH SEDATIVE, HYPNOTIC, OR ANXIOLYTIC-INDUCED DEPRESSIVE DISORDER
C0002726|T047|E85.9|DMDICD10|AMYLOIDOSIS, UNSPECIFIED|AMYLOIDOSE, NICHT NAEHER BEZEICHNET
C2878456|T037|T43.3X2A|ICD10CM|POISONING BY PHENOTHIAZINE ANTIPSYCHOTICS AND NEUROLEPTICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY PHENOTHIAZ ANTIPSYCHOT/NEUROLEPT, SELF-HARM, INIT
C2878458|T037|T43.3X2S|ICD10CM|POISONING BY PHENOTHIAZINE ANTIPSYCHOTICS AND NEUROLEPTICS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY PHENOTHIAZ ANTIPSYCHOT/NEUROLEPT, SLF-HRM, SEQUELA
C2893653|T047|M12.079|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], UNSPECIFIED ANKLE AND FOOT|CHRONIC POSTRHEUMATIC ARTHROPATHY, UNSP ANKLE AND FOOT
C3263952|T048|F03.91|ICD10CM|UNSPECIFIED DEMENTIA WITH BEHAVIORAL DISTURBANCE|UNSPECIFIED DEMENTIA WITH VIOLENT BEHAVIOR
C2833894|T037|S14.114A|ICD10CM|COMPLETE LESION AT C4 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION AT C4 LEVEL OF CERVICAL SPINAL CORD, INIT
C2882593|T047|I69.361|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING CEREBRAL INFARCTION AFFECTING RIGHT DOMINANT SIDE|OTH PARLYT SYNDROME FOL CEREB INFRC AFF RIGHT DOMINANT SIDE
C2882595|T047|I69.363|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING CEREBRAL INFARCTION AFFECTING RIGHT NON-DOMINANT SIDE|OTH PARLYT SYNDROME FOL CEREBRAL INFRC AFF RIGHT NONDOM SIDE
C2882594|T047|I69.362|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING CEREBRAL INFARCTION AFFECTING LEFT DOMINANT SIDE|OTH PARLYT SYNDROME FOL CEREB INFRC AFF LEFT DOMINANT SIDE
C2882597|T047|I69.365|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING CEREBRAL INFARCTION, BILATERAL|OTH PARALYTIC SYNDROME FOLLOWING CEREBRAL INFRC, BILATERAL
C2882596|T047|I69.364|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING CEREBRAL INFARCTION AFFECTING LEFT NON-DOMINANT SIDE|OTH PARLYT SYNDROME FOL CEREBRAL INFRC AFF LEFT NONDOM SIDE
C2882598|T047|I69.369|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING CEREBRAL INFARCTION AFFECTING UNSPECIFIED SIDE|OTH PARALYTIC SYNDROME FOL CEREBRAL INFRC AFF UNSP SIDE
C2891321|T037|T87.1X1|ICD10CM|COMPLICATIONS OF REATTACHED (PART OF) RIGHT LOWER EXTREMITY|COMPLICATIONS OF REATTACHED (PART OF) RIGHT LOWER EXTREMITY
C2860134|T037|S79.109A|ICD10CM|UNSPECIFIED PHYSEAL FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP PHYSEAL FRACTURE OF LOWER END OF UNSP FEMUR, INIT
C2842027|T191|C46.52|ICD10CM|KAPOSI'S SARCOMA OF LEFT LUNG|KAPOSI'S SARCOMA OF LEFT LUNG
C2842026|T191|C46.51|ICD10CM|KAPOSI'S SARCOMA OF RIGHT LUNG|KAPOSI'S SARCOMA OF RIGHT LUNG
C2888815|T047|M00.059|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, UNSPECIFIED HIP|STAPHYLOCOCCAL ARTHRITIS, UNSPECIFIED HIP
C2888814|T047|M00.052|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, LEFT HIP|STAPHYLOCOCCAL ARTHRITIS, LEFT HIP
C2888813|T047|M00.051|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, RIGHT HIP|STAPHYLOCOCCAL ARTHRITIS, RIGHT HIP
C2855842|T037|S68.012S|ICD10CM|COMPLETE TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF LEFT THUMB, SEQUELA|COMPLETE TRAUMATIC MCP AMPUTATION OF LEFT THUMB, SEQUELA
C2977711|T037|S02.609B|ICD10CM|FRACTURE OF MANDIBLE, UNSPECIFIED, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF MANDIBLE, UNSP, INIT ENCNTR FOR OPEN FRACTURE
C2977710|T037|S02.609A|ICD10CM|FRACTURE OF MANDIBLE, UNSPECIFIED, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF MANDIBLE, UNSP, INIT ENCNTR FOR CLOSED FRACTURE
C4270260|T046|T83.122A|ICD10CM|DISPLACEMENT OF INDWELLING URETERAL STENT, INITIAL ENCOUNTER|DISPLACEMENT OF INDWELLING URETERAL STENT, INITIAL ENCOUNTER
C2833622|T037|S12.650B|ICD10CM|OTHER TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH TRAUM DISPL SPONDYLOLYSIS OF 7TH CERVCAL VERT, 7THB
C0477976|T019|Q07.8|DMDICD10|OTHER SPECIFIED CONGENITAL MALFORMATIONS OF NERVOUS SYSTEM|SONSTIGE NAEHER BEZEICHNETE ANGEBORENE FEHLBILDUNGEN DES NERVENSYSTEMS
C2910110|T019|Q07.9|ICD10CM|CONGENITAL MALFORMATION OF NERVOUS SYSTEM, UNSPECIFIED|CONGENITAL DISEASE OR LESION NOS OF NERVOUS SYSTEM
C2885029|T037|T60.1X2S|ICD10CM|TOXIC EFFECT OF HALOGENATED INSECTICIDES, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF HALOGENATED INSECTICIDES, SELF-HARM, SEQUELA
C2977066|T047|J96.02|ICD10CM|ACUTE RESPIRATORY FAILURE WITH HYPERCAPNIA|ACUTE RESPIRATORY FAILURE WITH HYPERCAPNIA
C2977064|T047|J96.00|ICD10CM|ACUTE RESPIRATORY FAILURE, UNSPECIFIED WHETHER WITH HYPOXIA OR HYPERCAPNIA|ACUTE RESPIRATORY FAILURE, UNSP W HYPOXIA OR HYPERCAPNIA
C2977065|T047|J96.01|ICD10CM|ACUTE RESPIRATORY FAILURE WITH HYPOXIA|ACUTE RESPIRATORY FAILURE WITH HYPOXIA
C0348499|T047|E85.8|ICD10CM|OTHER AMYLOIDOSIS|OTHER AMYLOIDOSIS
C2874711|T048|F16.92|ICD10CM|HALLUCINOGEN USE, UNSPECIFIED WITH INTOXICATION, UNSPECIFIED|HALLUCINOGEN USE, UNSPECIFIED WITH INTOXICATION
C2874520|T048|F13.15|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED PSYCHOTIC DISORDER
C4509023|T047|E85.81|ICD10CM|LIGHT CHAIN (AL) AMYLOIDOSIS|LIGHT CHAIN (AL) AMYLOIDOSIS
C4237548|T048|F16.921|ICD10CM|HALLUCINOGEN USE, UNSPECIFIED WITH INTOXICATION WITH DELIRIUM|OTHER HALLUCINOGEN INTOXICATION DELIRIUM
C2874518|T048|F13.150|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|SEDATV/HYP/ANXIOLYTC ABUSE W PSYCHOTIC DISORDER W DELUSIONS
C4509024|T047|E85.82|ICD10CM|WILD-TYPE TRANSTHYRETIN-RELATED (ATTR) AMYLOIDOSIS|SENILE SYSTEMIC AMYLOIDOSIS (SSA)
C2833213|T037|S12.100B|ICD10CM|UNSPECIFIED DISPLACED FRACTURE OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP DISP FX OF SECOND CERVICAL VERTEBRA, INIT FOR OPN FX
C2833212|T037|S12.100A|ICD10CM|UNSPECIFIED DISPLACED FRACTURE OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP DISP FX OF SECOND CERVICAL VERTEBRA, INIT FOR CLOS FX
C2842138|T191|C50.919|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF UNSPECIFIED FEMALE BREAST|MALIGNANT NEOPLASM OF UNSP SITE OF UNSPECIFIED FEMALE BREAST
C2855859|T037|S68.029S|ICD10CM|PARTIAL TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF UNSPECIFIED THUMB, SEQUELA|PARTIAL TRAUMATIC MCP AMPUTATION OF THMB, SEQUELA
C0153687|T191|C79.2|DMDICD10|SECONDARY MALIGNANT NEOPLASM OF SKIN|SEKUNDAERE BOESARTIGE NEUBILDUNG DER HAUT
C2842136|T191|C50.911|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF RIGHT FEMALE BREAST|MALIGNANT NEOPLASM OF UNSP SITE OF RIGHT FEMALE BREAST
C2842137|T191|C50.912|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF LEFT FEMALE BREAST|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF LEFT FEMALE BREAST
C0036351|T048|F20.5|DMDICD10|RESIDUAL SCHIZOPHRENIA|SCHIZOPHRENES RESIDUUM
C2884721|T037|T57.92XA|ICD10CM|TOXIC EFFECT OF UNSPECIFIED INORGANIC SUBSTANCE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF UNSP INORGANIC SUBSTANCE, SELF-HARM, INIT
C0036349|T048|F20.0|DMDICD10|PARANOID SCHIZOPHRENIA|PARANOIDE SCHIZOPHRENIE
C0036347|T048|F20.1|DMDICD10|DISORGANIZED SCHIZOPHRENIA|HEBEPHRENE SCHIZOPHRENIE
C0036344|T048|F20.2|DMDICD10|CATATONIC SCHIZOPHRENIA|KATATONE SCHIZOPHRENIE
C0392322|T048|F20.3|DMDICD10|UNDIFFERENTIATED SCHIZOPHRENIA|UNDIFFERENZIERTE SCHIZOPHRENIE
C0036341|T048|F20.9|DMDICD10|SCHIZOPHRENIA, UNSPECIFIED|SCHIZOPHRENIE, NICHT NAEHER BEZEICHNET
C2859167|T037|S73.012A|ICD10CM|POSTERIOR SUBLUXATION OF LEFT HIP, INITIAL ENCOUNTER|POSTERIOR SUBLUXATION OF LEFT HIP, INITIAL ENCOUNTER
C2901798|T047|M86.121|ICD10CM|OTHER ACUTE OSTEOMYELITIS, RIGHT HUMERUS|OTHER ACUTE OSTEOMYELITIS, RIGHT HUMERUS
C2901799|T047|M86.122|ICD10CM|OTHER ACUTE OSTEOMYELITIS, LEFT HUMERUS|OTHER ACUTE OSTEOMYELITIS, LEFT HUMERUS
C2874163|T047|E13.610|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC NEUROPATHIC ARTHROPATHY|OTH DIABETES MELLITUS WITH DIABETIC NEUROPATHIC ARTHROPATHY
C2901800|T047|M86.129|ICD10CM|OTHER ACUTE OSTEOMYELITIS, UNSPECIFIED HUMERUS|OTHER ACUTE OSTEOMYELITIS, UNSPECIFIED HUMERUS
C2833998|T037|S14.142D|ICD10CM|BROWN-SEQUARD SYNDROME AT C2 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|BROWN-SEQUARD SYNDROME AT C2, SUBS
C2874164|T047|E13.618|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH OTHER DIABETIC ARTHROPATHY|OTH DIABETES MELLITUS WITH OTHER DIABETIC ARTHROPATHY
C2833997|T037|S14.142A|ICD10CM|BROWN-SEQUARD SYNDROME AT C2 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|BROWN-SEQUARD SYNDROME AT C2, INIT
C0349028|T191|D03.0|DMDICD10|MELANOMA IN SITU OF LIP|MELANOMA IN SITU DER LIPPE
C0349031|T191|D03.4|DMDICD10|MELANOMA IN SITU OF SCALP AND NECK|MELANOMA IN SITU DER BEHAARTEN KOPFHAUT UND DES HALSES
C0346040|T191|D03|DMDICD10|MELANOMA IN SITU, UNSPECIFIED|MELANOMA IN SITU
C1403733|T191||ICD10CM|MELANOMA IN SITU OF OTHER SITES
C2832134|T037|S06.319S|ICD10CM|CONTUSION AND LACERATION OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|CONTUS/LAC RIGHT CEREBRUM W LOC OF UNSP DURATION, SEQUELA
C2889289|T047|M05.569|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP KNEE
C2889287|T047|M05.561|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT KNEE|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889288|T047|M05.562|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT KNEE|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF LEFT KNEE
C0029640|T047|K56.4|ICD10CM|OTHER IMPACTION OF INTESTINE|OTHER IMPACTION OF INTESTINE
C0015734|T033||ICD10CM|FECAL IMPACTION
C2905701|T037|X74.01XS|ICD10CM|INTENTIONAL SELF-HARM BY AIRGUN, SEQUELA|INTENTIONAL SELF-HARM BY AIRGUN, SEQUELA
C2889262|T047|M05.49|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF MULTIPLE SITES
C2890830|T037|T84.610A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL FIXATION DEVICE OF RIGHT HUMERUS, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INT FIX OF RIGHT HUMERUS, INIT
C2889231|T047|M05.40|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSP SITE
C2905700|T037|X74.01XD|ICD10CM|INTENTIONAL SELF-HARM BY AIRGUN, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY AIRGUN, SUBSEQUENT ENCOUNTER
C2905699|T037|X74.01XA|ICD10CM|INTENTIONAL SELF-HARM BY AIRGUN, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY AIRGUN, INITIAL ENCOUNTER
C2905716|T037|X74.9XXA|ICD10CM|INTENTIONAL SELF-HARM BY UNSPECIFIED FIREARM DISCHARGE, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY UNSP FIREARM DISCHARGE, INIT ENCNTR
C2879390|T037|T46.0X2S|ICD10CM|POISONING BY CARDIAC-STIMULANT GLYCOSIDES AND DRUGS OF SIMILAR ACTION, INTENTIONAL SELF-HARM, SEQUELA|POISN BY CARDI-STIM GLYCOS/DRUG SIMLAR ACT, SLF-HRM, SEQUELA
C2905717|T037|X74.9XXD|ICD10CM|INTENTIONAL SELF-HARM BY UNSPECIFIED FIREARM DISCHARGE, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY UNSP FIREARM DISCHARGE, SUBS ENCNTR
C2905718|T037|X74.9XXS|ICD10CM|INTENTIONAL SELF-HARM BY UNSPECIFIED FIREARM DISCHARGE, SEQUELA|INTENTIONAL SELF-HARM BY UNSP FIREARM DISCHARGE, SEQUELA
C2856896|T037|S72.051A|ICD10CM|UNSPECIFIED FRACTURE OF HEAD OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF HEAD OF RIGHT FEMUR, INIT FOR CLOS FX
C2856898|T037|S72.051C|ICD10CM|UNSPECIFIED FRACTURE OF HEAD OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP FX HEAD OF RIGHT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2856897|T037|S72.051B|ICD10CM|UNSPECIFIED FRACTURE OF HEAD OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP FX HEAD OF RIGHT FEMUR, INIT FOR OPN FX TYPE I/2
C2901553|T046|M84.672A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, LEFT ANKLE, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, LEFT ANKLE, INIT
C2900548|T046|M80.871A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, RIGHT ANKLE AND FOOT, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, RIGHT ANK/FT, INIT
C2838437|T037|S32.612B|ICD10CM|DISPLACED AVULSION FRACTURE OF LEFT ISCHIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISPLACED AVULSION FRACTURE OF LEFT ISCHIUM, INIT FOR OPN FX
C2838436|T037|S32.612A|ICD10CM|DISPLACED AVULSION FRACTURE OF LEFT ISCHIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED AVULSION FRACTURE OF LEFT ISCHIUM, INIT
C2837617|T037|S32.049A|ICD10CM|UNSPECIFIED FRACTURE OF FOURTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF FOURTH LUMBAR VERTEBRA, INIT FOR CLOS FX
C0564750|T046||ICD10CM|EMBOLISM AND THROMBOSIS OF ARTERIES OF EXTREMITIES, UNSPECIFIED
C0155755|T046|I74.5|DMDICD10|EMBOLISM AND THROMBOSIS OF ILIAC ARTERY|EMBOLIE UND THROMBOSE DER A. ILIACA
C4270256|T046|T83.113A|ICD10CM|BREAKDOWN (MECHANICAL) OF OTHER URINARY STENTS, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF OTHER URINARY STENTS, INIT
C2837618|T037|S32.049B|ICD10CM|UNSPECIFIED FRACTURE OF FOURTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF FOURTH LUMBAR VERTEBRA, INIT FOR OPN FX
C0494620|T046|I74.2|DMDICD10|EMBOLISM AND THROMBOSIS OF ARTERIES OF THE UPPER EXTREMITIES|EMBOLIE UND THROMBOSE DER ARTERIEN DER OBEREN EXTREMITAETEN
C0340589|T046|I74.3|DMDICD10|EMBOLISM AND THROMBOSIS OF ARTERIES OF THE LOWER EXTREMITIES|EMBOLIE UND THROMBOSE DER ARTERIEN DER UNTEREN EXTREMITAETEN
C0348650|T047|I74.8|DMDICD10|EMBOLISM AND THROMBOSIS OF OTHER ARTERIES|EMBOLIE UND THROMBOSE SONSTIGER ARTERIEN
C0013924|T046|I74.9|DMDICD10|EMBOLISM AND THROMBOSIS OF UNSPECIFIED ARTERY|EMBOLIE UND THROMBOSE NICHT NAEHER BEZEICHNETER ARTERIE
C2900961|T046|M84.443A|ICD10CM|PATHOLOGICAL FRACTURE, UNSPECIFIED HAND, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, UNSP HAND, INIT ENCNTR FOR FRACTURE
C2901466|T046|M84.649A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, UNSPECIFIED HAND, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, UNSP HAND, INIT FOR FX
C2833317|T037|S12.200B|ICD10CM|UNSPECIFIED DISPLACED FRACTURE OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP DISP FX OF THIRD CERVICAL VERTEBRA, INIT FOR OPN FX
C2833316|T037|S12.200A|ICD10CM|UNSPECIFIED DISPLACED FRACTURE OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP DISP FX OF THIRD CERVICAL VERTEBRA, INIT FOR CLOS FX
C0839952|T047|M86.249|ICD10CM|SUBACUTE OSTEOMYELITIS, UNSPECIFIED HAND|SUBACUTE OSTEOMYELITIS, UNSPECIFIED HAND
C4268058|T047|E10.3559|ICD10CM|TYPE 1 DIABETES MELLITUS WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, UNSPECIFIED EYE|TYPE 1 DIABETES WITH STABLE PROLIF DIABETIC RTNOP, UNSP
C4268056|T047|E10.3552|ICD10CM|TYPE 1 DIABETES MELLITUS WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, LEFT EYE|TYPE 1 DIABETES WITH STABLE PROLIF DIABETIC RTNOP, LEFT EYE
C4268057|T047|E10.3553|ICD10CM|TYPE 1 DIABETES MELLITUS WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, BILATERAL|TYPE 1 DIABETES WITH STABLE PROLIF DIABETIC RTNOP, BILATERAL
C4268055|T047|E10.3551|ICD10CM|TYPE 1 DIABETES MELLITUS WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, RIGHT EYE|TYPE 1 DIABETES WITH STABLE PROLIF DIABETIC RTNOP, RIGHT EYE
C2858852|T037|S72.461B|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL SUPRCNDL FX W INTRCNDL EXTN LOW END R FEMR, 7THB
C2858853|T037|S72.461C|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL SUPRCNDL FX W INTRCNDL EXTN LOW END R FEMR, 7THC
C2834036|T037|S14.152A|ICD10CM|OTHER INCOMPLETE LESION AT C2 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|OTH INCOMPLETE LESION AT C2, INIT
C4268241|T048|F14.94|ICD10CM|COCAINE USE, UNSPECIFIED WITH COCAINE-INDUCED MOOD DISORDER|COCAINE INDUCED BIPOLAR OR RELATED DISORDER, WITHOUT USE DISORDER
C2858593|T037|S72.434A|ICD10CM|NONDISPLACED FRACTURE OF MEDIAL CONDYLE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF MEDIAL CONDYLE OF RIGHT FEMUR, INIT
C2882743|T047|I70.299|ICD10CM|OTHER ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES, UNSPECIFIED EXTREMITY|OTH ATHSCL NATIVE ARTERIES OF EXTREMITIES, UNSP EXTREMITY
C2882742|T047|I70.298|ICD10CM|OTHER ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES, OTHER EXTREMITY|OTH ATHSCL NATIVE ARTERIES OF EXTREMITIES, OTH EXTREMITY
C3264138|T033|Z89.519|ICD10CM|ACQUIRED ABSENCE OF UNSPECIFIED LEG BELOW KNEE|ACQUIRED ABSENCE OF UNSPECIFIED LEG BELOW KNEE
C2882741|T047|I70.293|ICD10CM|OTHER ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES, BILATERAL LEGS|OTH ATHSCL NATIVE ARTERIES OF EXTREMITIES, BILATERAL LEGS
C2882740|T047|I70.292|ICD10CM|OTHER ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES, LEFT LEG|OTH ATHSCL NATIVE ARTERIES OF EXTREMITIES, LEFT LEG
C2882739|T047|I70.291|ICD10CM|OTHER ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES, RIGHT LEG|OTH ATHSCL NATIVE ARTERIES OF EXTREMITIES, RIGHT LEG
C2834038|T037|S14.152S|ICD10CM|OTHER INCOMPLETE LESION AT C2 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|OTH INCOMPLETE LESION AT C2, SEQUELA
C2905752|T037|X78.0XXS|ICD10CM|INTENTIONAL SELF-HARM BY SHARP GLASS, SEQUELA|INTENTIONAL SELF-HARM BY SHARP GLASS, SEQUELA
C2832284|T037|S06.355S|ICD10CM|TRAUMATIC HEMORRHAGE OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, SEQUELA|TRAUM HEMOR L CEREB W LOC >24 HR W RET CONSC LEV, SEQUELA
C2890731|T037|T84.290A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTERNAL FIXATION DEVICE OF BONES OF HAND AND FINGERS, INITIAL ENCOUNTER|MECH COMPL OF INT FIX OF BONES OF HAND AND FINGERS, INIT
C2832076|T037|S06.305S|ICD10CM|UNSPECIFIED FOCAL TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, SEQUELA|UNSP FOCAL TBI W LOC >24 HR W RET CONSC LEV, SEQUELA
C2887458|T047||ICD10CM|MODERATE PERSISTENT ASTHMA WITH STATUS ASTHMATICUS
C2887456|T047||ICD10CM|MODERATE PERSISTENT ASTHMA, UNCOMPLICATED
C2887457|T033||ICD10CM|MODERATE PERSISTENT ASTHMA WITH (ACUTE) EXACERBATION
C2832074|T037|S06.305A|ICD10CM|UNSPECIFIED FOCAL TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, INITIAL ENCOUNTER|UNSP FOCAL TBI W LOC >24 HR W RET CONSC LEV, INIT
C2883012|T047|I70.749|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF UNSPECIFIED SITE|ATHSCL TYPE OF BYPASS OF THE LEFT LEG W ULCER OF UNSP SITE
C2883011|T047|I70.748|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF OTHER PART OF LOWER LEG|ATHSCL TYPE OF BYPASS OF LEFT LEG W ULCER OTH PRT LOW LEG
C2883004|T047|I70.741|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF THIGH|ATHSCL TYPE OF BYPASS OF THE LEFT LEG W ULCERATION OF THIGH
C4269245|T037|S02.109B|ICD10CM|FRACTURE OF BASE OF SKULL, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF BASE OF SKULL, UNSPECIFIED SIDE, 7THB
C2883006|T047|I70.743|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF ANKLE|ATHSCL TYPE OF BYPASS OF THE LEFT LEG W ULCERATION OF ANKLE
C2883005|T047|I70.742|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF CALF|ATHSCL TYPE OF BYPASS OF THE LEFT LEG W ULCERATION OF CALF
C2883010|T047|I70.745|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF OTHER PART OF FOOT|ATHSCL TYPE OF BYPASS OF THE LEFT LEG W ULCER OTH PRT FOOT
C2883008|T047|I70.744|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF HEEL AND MIDFOOT|ATHSCL TYPE OF BYPASS OF LEFT LEG W ULCER OF HEEL AND MIDFT
C4269494|T037|S02.631S|ICD10CM|FRACTURE OF CORONOID PROCESS OF RIGHT MANDIBLE, SEQUELA|FRACTURE OF CORONOID PROCESS OF RIGHT MANDIBLE, SEQUELA
C2874577|T048||ICD10CM|COCAINE ABUSE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE
C2888919|T047|M00.869|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, UNSPECIFIED KNEE|ARTHRITIS DUE TO OTHER BACTERIA, UNSPECIFIED KNEE
C2874576|T048|F14.121|ICD10CM|COCAINE ABUSE WITH INTOXICATION WITH DELIRIUM|COCAINE ABUSE WITH INTOXICATION WITH DELIRIUM
C2888918|T047|M00.862|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, LEFT KNEE|ARTHRITIS DUE TO OTHER BACTERIA, LEFT KNEE
C2888917|T047|M00.861|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, RIGHT KNEE|ARTHRITIS DUE TO OTHER BACTERIA, RIGHT KNEE
C2874578|T048|F14.129|ICD10CM|COCAINE ABUSE WITH INTOXICATION, UNSPECIFIED|COCAINE ABUSE WITH INTOXICATION, UNSPECIFIED
C2888234|T047|L89.009|ICD10CM|PRESSURE ULCER OF UNSPECIFIED ELBOW, UNSPECIFIED STAGE|HEALING PRESSURE ULCER OF UNSPECIFIED ELBOW, UNSPECIFIED STAGE
C2888207|T047|L89.001|ICD10CM|PRESSURE ULCER OF UNSPECIFIED ELBOW, STAGE 1|PRESSURE ULCER OF UNSPECIFIED ELBOW, STAGE 1
C2888204|T047|L89.000|ICD10CM|PRESSURE ULCER OF UNSPECIFIED ELBOW, UNSTAGEABLE|PRESSURE ULCER OF UNSPECIFIED ELBOW, UNSTAGEABLE
C2888213|T047|L89.003|ICD10CM|PRESSURE ULCER OF UNSPECIFIED ELBOW, STAGE 3|PRESSURE ULCER OF UNSPECIFIED ELBOW, STAGE 3
C2888210|T047|L89.002|ICD10CM|PRESSURE ULCER OF UNSPECIFIED ELBOW, STAGE 2|PRESSURE ULCER OF UNSPECIFIED ELBOW, STAGE 2
C2888216|T047|L89.004|ICD10CM|PRESSURE ULCER OF UNSPECIFIED ELBOW, STAGE 4|PRESSURE ULCER OF UNSPECIFIED ELBOW, STAGE 4
C2857873|T037|S72.334A|ICD10CM|NONDISPLACED OBLIQUE FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED OBLIQUE FRACTURE OF SHAFT OF RIGHT FEMUR, INIT
C2857875|T037|S72.334C|ICD10CM|NONDISPLACED OBLIQUE FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP OBLIQUE FX SHAFT OF R FEMR, 7THC
C2857874|T037|S72.334B|ICD10CM|NONDISPLACED OBLIQUE FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP OBLIQUE FX SHAFT OF R FEMR, INIT FOR OPN FX TYPE I/2
C2882919|T047|I70.608|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, OTHER EXTREMITY|UNSP ATHSCL NONBIOL BYPASS OF THE EXTREMITIES, OTH EXTREMITY
C2882920|T047|I70.609|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, UNSPECIFIED EXTREMITY|UNSP ATHSCL NONBIOL BYPASS OF THE EXTRM, UNSP EXTREMITY
C2882916|T047|I70.601|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, RIGHT LEG|UNSP ATHSCL NONBIOL BYPASS OF THE EXTREMITIES, RIGHT LEG
C2882917|T047|I70.602|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, LEFT LEG|UNSP ATHSCL NONBIOL BYPASS OF THE EXTREMITIES, LEFT LEG
C2882918|T047|I70.603|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, BILATERAL LEGS|UNSP ATHSCL NONBIOL BYPASS OF THE EXTRM, BILATERAL LEGS
C2901937|T046|M87.011|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF RIGHT SHOULDER|IDIOPATHIC ASEPTIC NECROSIS OF RIGHT SHOULDER
C2860023|T037|S78.911A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT HIP AND THIGH, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMP OF R HIP AND THIGH, LEVEL UNSP, INIT
C2860075|T037|S79.011A|ICD10CM|SALTER-HARRIS TYPE I PHYSEAL FRACTURE OF UPPER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SLTR-HARIS TYPE I PHYSEAL FX UPPER END OF RIGHT FEMUR, INIT
C2860024|T037|S78.911D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT HIP AND THIGH, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMP OF R HIP AND THIGH, LEVEL UNSP, SUBS
C2890658|T037|T84.190A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTERNAL FIXATION DEVICE OF RIGHT HUMERUS, INITIAL ENCOUNTER|MECH COMPL OF INT FIX OF RIGHT HUMERUS, INIT
C0266460|T019||ICD10CM|MICROCEPHALY
C2837502|T037|S32.018A|ICD10CM|OTHER FRACTURE OF FIRST LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF FIRST LUMBAR VERTEBRA, INIT FOR CLOS FX
C2832527|T037|S06.6X4S|ICD10CM|TRAUMATIC SUBARACHNOID HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|TRAUM SUBRAC HEM W LOC OF 6 HOURS TO 24 HOURS, SEQUELA
C2901886|T047|M86.469|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, UNSPECIFIED TIBIA AND FIBULA|CHRONIC OSTEOMYELIT W DRAINING SINUS, UNSP TIBIA AND FIBULA
C2869770|T037|S98.021S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT FOOT AT ANKLE LEVEL, SEQUELA|PARTIAL TRAUMATIC AMP OF RIGHT FOOT AT ANKLE LEVEL, SEQUELA
C2885141|T037|T61.12XS|ICD10CM|SCOMBROID FISH POISONING, INTENTIONAL SELF-HARM, SEQUELA|SCOMBROID FISH POISONING, INTENTIONAL SELF-HARM, SEQUELA
C2901884|T047|M86.461|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, RIGHT TIBIA AND FIBULA|CHRONIC OSTEOMYELIT W DRAINING SINUS, RIGHT TIBIA AND FIBULA
C2901885|T047|M86.462|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, LEFT TIBIA AND FIBULA|CHRONIC OSTEOMYELIT W DRAINING SINUS, LEFT TIBIA AND FIBULA
C2885139|T037|T61.12XA|ICD10CM|SCOMBROID FISH POISONING, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|SCOMBROID FISH POISONING, INTENTIONAL SELF-HARM, INIT ENCNTR
C2869768|T037|S98.021A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT FOOT AT ANKLE LEVEL, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP OF RIGHT FOOT AT ANKLE LEVEL, INIT
C2869769|T037|S98.021D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT FOOT AT ANKLE LEVEL, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMP OF RIGHT FOOT AT ANKLE LEVEL, SUBS
C2832236|T037|S06.344A|ICD10CM|TRAUMATIC HEMORRHAGE OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|TRAUM HEMOR RIGHT CEREBRUM W LOC OF 6-24 HRS, INIT
C2884578|T037|T56.7X2S|ICD10CM|TOXIC EFFECT OF BERYLLIUM AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF BERYLLIUM AND ITS COMPND, SELF-HARM, SEQUELA
C2859256|T037|S73.046A|ICD10CM|CENTRAL DISLOCATION OF UNSPECIFIED HIP, INITIAL ENCOUNTER|CENTRAL DISLOCATION OF UNSPECIFIED HIP, INITIAL ENCOUNTER
C2832238|T037|S06.344S|ICD10CM|TRAUMATIC HEMORRHAGE OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|TRAUM HEMOR RIGHT CEREBRUM W LOC OF 6-24 HRS, SEQUELA
C2874775|T048|F18.920|ICD10CM|INHALANT USE, UNSPECIFIED WITH INTOXICATION, UNCOMPLICATED|INHALANT USE, UNSPECIFIED WITH INTOXICATION, UNCOMPLICATED
C2874776|T048|F18.921|ICD10CM|INHALANT USE, UNSPECIFIED WITH INTOXICATION WITH DELIRIUM|INHALANT USE, UNSPECIFIED WITH INTOXICATION WITH DELIRIUM
C2869803|T037|S98.129D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED GREAT TOE, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF UNSP GREAT TOE, SUBS ENCNTR
C2884576|T037|T56.7X2A|ICD10CM|TOXIC EFFECT OF BERYLLIUM AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF BERYLLIUM AND ITS COMPOUNDS, SELF-HARM, INIT
C2874219|T047|E44.1|ICD10CM|MILD PROTEIN-CALORIE MALNUTRITION|MILD PROTEIN-CALORIE MALNUTRITION
C2874777|T048|F18.929|ICD10CM|INHALANT USE, UNSPECIFIED WITH INTOXICATION, UNSPECIFIED|INHALANT USE, UNSPECIFIED WITH INTOXICATION, UNSPECIFIED
C2861639|T191||ICD10CM|ACUTE PANMYELOSIS WITH MYELOFIBROSIS, IN REMISSION
C2861638|T191|C94.40|ICD10CM|ACUTE PANMYELOSIS WITH MYELOFIBROSIS NOT HAVING ACHIEVED REMISSION|ACUTE PANMYELOSIS W MYELOFIBROSIS NOT ACHIEVE REMISSION
C2861640|T191||ICD10CM|ACUTE PANMYELOSIS WITH MYELOFIBROSIS, IN RELAPSE
C2883076|T047|I80.291|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF OTHER DEEP VESSELS OF RIGHT LOWER EXTREMITY|PHLEBITIS AND THOMBOPHLB OF DEEP VESSELS OF R LOW EXTREM
C2883077|T047|I80.292|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF OTHER DEEP VESSELS OF LEFT LOWER EXTREMITY|PHLEBITIS AND THOMBOPHLB OF DEEP VESSELS OF L LOW EXTREM
C2883078|T047|I80.293|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF OTHER DEEP VESSELS OF LOWER EXTREMITY, BILATERAL|PHLEBITIS AND THOMBOPHLB OF DEEP VESSELS OF LOW EXTRM, BI
C2883079|T047|I80.299|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF OTHER DEEP VESSELS OF UNSPECIFIED LOWER EXTREMITY|PHLEBITIS AND THOMBOPHLB OF DEEP VESSELS OF UNSP LOW EXTRM
C2874013|T047|E09.69|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATION|DRUG/CHEM DIABETES MELLITUS W OTH COMPLICATION
C2874749|T048|F18.129|ICD10CM|INHALANT ABUSE WITH INTOXICATION, UNSPECIFIED|INHALANT ABUSE WITH INTOXICATION, UNSPECIFIED
C2874012|T047|E09.65|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH HYPERGLYCEMIA|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS W HYPERGLYCEMIA
C2878947|T037|T44.8X2A|ICD10CM|POISONING BY CENTRALLY-ACTING AND ADRENERGIC-NEURON-BLOCKING AGENTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY CENTR-ACTING/ADREN-NEURN-BLOCK AGNT, SLF-HRM, INIT
C2877122|T037|T38.5X2A|ICD10CM|POISONING BY OTHER ESTROGENS AND PROGESTOGENS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH ESTROGENS AND PROGESTOGENS, SELF-HARM, INIT
C2874896|T048|F31.64|ICD10CM|BIPOLAR DISORDER, CURRENT EPISODE MIXED, SEVERE, WITH PSYCHOTIC FEATURES|BIPOLAR DISORD, CRNT EPISODE MIXED, SEVERE, W PSYCH FEATURES
C2874891|T048|F31.61|ICD10CM|BIPOLAR DISORDER, CURRENT EPISODE MIXED, MILD|BIPOLAR DISORDER, CURRENT EPISODE MIXED, MILD
C2874890|T048|F31.6|ICD10CM|BIPOLAR DISORDER, CURRENT EPISODE MIXED, UNSPECIFIED|BIPOLAR DISORDER, CURRENT EPISODE MIXED
C2874893|T048|F31.63|ICD10CM|BIPOLAR DISORDER, CURRENT EPISODE MIXED, SEVERE, WITHOUT PSYCHOTIC FEATURES|BIPOLAR DISORD, CRNT EPSD MIXED, SEVERE, W/O PSYCH FEATURES
C2874892|T048|F31.62|ICD10CM|BIPOLAR DISORDER, CURRENT EPISODE MIXED, MODERATE|BIPOLAR DISORDER, CURRENT EPISODE MIXED, MODERATE
C2349274|T191|C91.92|ICD10CM|LYMPHOID LEUKEMIA, UNSPECIFIED, IN RELAPSE|LYMPHOID LEUKEMIA, UNSPECIFIED, IN RELAPSE
C0686597|T191||ICD10AM|LYMPHOID LEUKEMIA, UNSPECIFIED, IN REMISSION
C2854113|T191|C91.90|ICD10CM|LYMPHOID LEUKEMIA, UNSPECIFIED NOT HAVING ACHIEVED REMISSION|LYMPHOID LEUKEMIA, UNSPECIFIED NOT HAVING ACHIEVED REMISSION
C2838079|T037|S32.425B|ICD10CM|NONDISPLACED FRACTURE OF POSTERIOR WALL OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP FX OF POSTERIOR WALL OF LEFT ACETAB, INIT FOR OPN FX
C2838078|T037|S32.425A|ICD10CM|NONDISPLACED FRACTURE OF POSTERIOR WALL OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF POSTERIOR WALL OF LEFT ACETABULUM, INIT
C2874748|T048|F18.121|ICD10CM|INHALANT ABUSE WITH INTOXICATION DELIRIUM|INHALANT ABUSE WITH INTOXICATION DELIRIUM
C4268079|T047|E11.3319|ICD10CM|TYPE 2 DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|TYPE 2 DIAB WITH MOD NONP RTNOP WITH MACULAR EDEMA, UNSP
C2882295|T047|I60.11|ICD10CM|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM RIGHT MIDDLE CEREBRAL ARTERY|NTRM SUBARACH HEMORRHAGE FROM RIGHT MIDDLE CEREBRAL ARTERY
C2882294|T047|I60.10|ICD10CM|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM UNSPECIFIED MIDDLE CEREBRAL ARTERY|NTRM SUBARACH HEMORRHAGE FROM UNSP MIDDLE CEREBRAL ARTERY
C2882296|T047|I60.12|ICD10CM|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM LEFT MIDDLE CEREBRAL ARTERY|NTRM SUBARACH HEMORRHAGE FROM LEFT MIDDLE CEREBRAL ARTERY
C4268076|T047|E11.3311|ICD10CM|TYPE 2 DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|TYPE 2 DIAB WITH MOD NONP RTNOP WITH MACULAR EDEMA, R EYE
C4268078|T047|E11.3313|ICD10CM|TYPE 2 DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|TYPE 2 DIAB WITH MODERATE NONP RTNOP WITH MACULAR EDEMA, BI
C4268077|T047|E11.3312|ICD10CM|TYPE 2 DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|TYPE 2 DIAB WITH MOD NONP RTNOP WITH MACULAR EDEMA, L EYE
C2874255|T047|E71.548|ICD10CM|OTHER PEROXISOMAL DISORDERS|OTHER PEROXISOMAL DISORDERS
C4270419|T046|T83.729A|ICD10CM|EXPOSURE OF OTHER PROSTHETIC MATERIALS INTO ORGAN OR TISSUE, INITIAL ENCOUNTER|EXPOSURE OF OTHER PROSTH MATRL INTO ORGAN OR TISSUE, INIT
C0751552|T191|C37|DMDICD10|MALIGNANT NEOPLASM OF THYMUS|BOESARTIGE NEUBILDUNG DES THYMUS
C0282529|T047||ICD10CM|RHIZOMELIC CHONDRODYSPLASIA PUNCTATA
C0751594|T047||ICD10CM|ZELLWEGER-LIKE SYNDROME
C2874256|T047|E71.542|ICD10CM|OTHER GROUP 3 PEROXISOMAL DISORDERS|OTHER GROUP 3 PEROXISOMAL DISORDERS
C2832449|T037|S06.4X5A|ICD10CM|EPIDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, INITIAL ENCOUNTER|EPIDURAL HEMORRHAGE W LOC >24 HR W RET CONSC LEV, INIT
C2879493|T037|T46.4X2S|ICD10CM|POISONING BY ANGIOTENSIN-CONVERTING-ENZYME INHIBITORS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY ANGIOTENS-CONVERT-ENZYME INHIBTR, SLF-HRM, SEQUELA
C2890284|T037|T83.191A|ICD10CM|OTHER MECHANICAL COMPLICATION OF IMPLANTED URINARY SPHINCTER, INITIAL ENCOUNTER|MECH COMPL OF IMPLANTED URINARY SPHINCTER, INITIAL ENCOUNTER
C2832451|T037|S06.4X5S|ICD10CM|EPIDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, SEQUELA|EPIDURAL HEMORRHAGE W LOC >24 HR W RET CONSC LEV, SEQUELA
C2877124|T037|T38.5X2S|ICD10CM|POISONING BY OTHER ESTROGENS AND PROGESTOGENS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH ESTROGENS AND PROGSTRN, SELF-HARM, SEQUELA
C2879491|T037|T46.4X2A|ICD10CM|POISONING BY ANGIOTENSIN-CONVERTING-ENZYME INHIBITORS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY ANGIOTENS-CONVERT-ENZYME INHIBTR, SELF-HARM, INIT
C2905680|T037|X73.1XXD|ICD10CM|INTENTIONAL SELF-HARM BY HUNTING RIFLE DISCHARGE, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY HUNTING RIFLE DISCHARGE, SUBS
C2902073|T046|M87.273|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED ANKLE|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED ANKLE
C2832175|T037|S06.329S|ICD10CM|CONTUSION AND LACERATION OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|CONTUS/LAC LEFT CEREBRUM W LOC OF UNSP DURATION, SEQUELA
C2875174|T047|G43.709|ICD10CM|CHRONIC MIGRAINE WITHOUT AURA, NOT INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|CHRONIC MIGRAINE W/O AURA, NOT INTRACTABLE, W/O STAT MIGR
C2901379|T046|M84.612A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, LEFT SHOULDER, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, LEFT SHOULDER, INIT
C2905758|T037|X78.2XXA|ICD10CM|INTENTIONAL SELF-HARM BY SWORD OR DAGGER, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY SWORD OR DAGGER, INITIAL ENCOUNTER
C2875173|T047|G43.701|ICD10CM|CHRONIC MIGRAINE WITHOUT AURA, NOT INTRACTABLE, WITH STATUS MIGRAINOSUS|CHRONIC MIGRAINE W/O AURA, NOT INTRACTABLE, W STAT MIGR
C2837660|T037|S32.10XA|ICD10CM|UNSPECIFIED FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF SACRUM, INIT ENCNTR FOR CLOSED FRACTURE
C2855915|T037|S68.122S|ICD10CM|PARTIAL TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF RIGHT MIDDLE FINGER, SEQUELA|PARTIAL TRAUMATIC MCP AMPUTATION OF R MID FINGER, SEQUELA
C2888883|T047|M00.261|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, RIGHT KNEE|OTHER STREPTOCOCCAL ARTHRITIS, RIGHT KNEE
C2859061|T037|S72.8X9A|ICD10CM|OTHER FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF UNSP FEMUR, INIT ENCNTR FOR CLOSED FRACTURE
C2859062|T037|S72.8X9B|ICD10CM|OTHER FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|OTH FRACTURE OF UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2888884|T047|M00.262|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, LEFT KNEE|OTHER STREPTOCOCCAL ARTHRITIS, LEFT KNEE
C2885713|T037|T63.482S|ICD10CM|TOXIC EFFECT OF VENOM OF OTHER ARTHROPOD, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF ARTHROPOD, SELF-HARM, SEQUELA
C2888885|T047|M00.269|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, UNSPECIFIED KNEE|OTHER STREPTOCOCCAL ARTHRITIS, UNSPECIFIED KNEE
C0013720|T047|Q79.6|DMDICD10|EHLERS-DANLOS SYNDROME|EHLERS-DANLOS-SYNDROM
C2857291|T037|S72.123A|ICD10CM|DISPLACED FRACTURE OF LESSER TROCHANTER OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF LESSER TROCHANTER OF UNSP FEMUR, INIT FOR CLOS FX
C2895335|T037|M48.56XA|ICD10CM|COLLAPSED VERTEBRA, NOT ELSEWHERE CLASSIFIED, LUMBAR REGION, INITIAL ENCOUNTER FOR FRACTURE|COLLAPSED VERTEBRA, NEC, LUMBAR REGION, INIT
C2883143|T047|I82.599|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF OTHER SPECIFIED DEEP VEIN OF UNSPECIFIED LOWER EXTREMITY|CHRONIC EMBOLISM AND THOMBOS OF DEEP VEIN OF UNSP LOW EXTRM
C0025269|T191|E31.23|ICD10CM|MULTIPLE ENDOCRINE NEOPLASIA [MEN] TYPE IIB|MULTIPLE ENDOCRINE NEOPLASIA [MEN] TYPE IIB
C0027662|T047|E31.20|ICD10CM|MULTIPLE ENDOCRINE NEOPLASIA [MEN] SYNDROME, UNSPECIFIED|MULTIPLE ENDOCRINE NEOPLASIA [MEN] SYNDROME, UNSPECIFIED
C0025267|T191|E31.21|ICD10CM|MULTIPLE ENDOCRINE NEOPLASIA [MEN] TYPE I|MULTIPLE ENDOCRINE NEOPLASIA [MEN] TYPE I
C2883140|T047|I82.591|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF OTHER SPECIFIED DEEP VEIN OF RIGHT LOWER EXTREMITY|CHRONIC EMBOLISM AND THROMBOSIS OF DEEP VEIN OF R LOW EXTREM
C2883142|T047|I82.593|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF OTHER SPECIFIED DEEP VEIN OF LOWER EXTREMITY, BILATERAL|CHRONIC EMBOLISM AND THOMBOS OF DEEP VEIN OF LOW EXTRM, BI
C2883141|T047|I82.592|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF OTHER SPECIFIED DEEP VEIN OF LEFT LOWER EXTREMITY|CHRONIC EMBOLISM AND THROMBOSIS OF DEEP VEIN OF L LOW EXTREM
C2832592|T037|S06.820S|ICD10CM|INJURY OF LEFT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|INJURY OF L INT CAROTID, INTCR W/O LOC, SEQUELA
C2910133|T019|Q24.5|ICD10CM|MALFORMATION OF CORONARY VESSELS|CONGENITAL CORONARY (ARTERY) ANEURYSM
C2837531|T037|S32.022A|ICD10CM|UNSTABLE BURST FRACTURE OF SECOND LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSTABLE BURST FRACTURE OF SECOND LUMBAR VERTEBRA, INIT
C2889544|T047|M08.06|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED KNEE|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, KNEE
C0155789|T047||ICD10CM|ESOPHAGEAL VARICES WITH BLEEDING
C0267092|T047|I85.00|ICD10CM|ESOPHAGEAL VARICES WITHOUT BLEEDING|ESOPHAGEAL VARICES WITHOUT BLEEDING
C2889543|T047|M08.062|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, LEFT KNEE|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, LEFT KNEE
C2889542|T047|M08.061|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, RIGHT KNEE|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, RIGHT KNEE
C4270585|T046|T85.733A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO IMPLANTED ELECTRONIC NEUROSTIMULATOR OF SPINAL CORD, ELECTRODE (LEAD), INITIAL ENCOUNTER|I/I REACT D/T IMPLNT ELEC NSTIM OF SPINAL CORD, LEAD, INIT
C2833880|T037|S14.109S|ICD10CM|UNSPECIFIED INJURY AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, SEQUELA|UNSP INJURY AT UNSP LEVEL OF CERVICAL SPINAL CORD, SEQUELA
C2832173|T037|S06.329A|ICD10CM|CONTUSION AND LACERATION OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|CONTUS/LAC LEFT CEREBRUM W LOC OF UNSP DURATION, INIT
C2885460|T037|T63.112S|ICD10CM|TOXIC EFFECT OF VENOM OF GILA MONSTER, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF GILA MONSTER, SELF-HARM, SEQUELA
C0837511|T047|M05.049|ICD10CM|FELTY'S SYNDROME, UNSPECIFIED HAND|FELTY'S SYNDROME, UNSPECIFIED HAND
C2889121|T047|M05.042|ICD10CM|FELTY'S SYNDROME, LEFT HAND|FELTY'S SYNDROME, LEFT HAND
C2889120|T047|M05.041|ICD10CM|FELTY'S SYNDROME, RIGHT HAND|FELTY'S SYNDROME, RIGHT HAND
C2887063|T047||ICD10CM|DIPHTHERITIC CARDIOMYOPATHY
C2887066|T047|A36.84|ICD10CM|DIPHTHERITIC TUBULO-INTERSTITIAL NEPHROPATHY|DIPHTHERITIC TUBULO-INTERSTITIAL NEPHROPATHY
C2902013|T046|M87.159|ICD10CM|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED FEMUR|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED FEMUR
C2902012|T046|M87.152|ICD10CM|OSTEONECROSIS DUE TO DRUGS, LEFT FEMUR|OSTEONECROSIS DUE TO DRUGS, LEFT FEMUR
C2902010|T047||ICD10CM|OSTEONECROSIS DUE TO DRUGS, PELVIS
C2902011|T046|M87.151|ICD10CM|OSTEONECROSIS DUE TO DRUGS, RIGHT FEMUR|OSTEONECROSIS DUE TO DRUGS, RIGHT FEMUR
C2910371|T047|Q93.88|ICD10CM|OTHER MICRODELETIONS|OTHER MICRODELETIONS
C0005138|T037|J63.2|DMDICD10|BERYLLIOSIS|BERYLLIOSE
C2853891|T191|C83.07|ICD10CM|SMALL CELL B-CELL LYMPHOMA, SPLEEN|SMALL CELL B-CELL LYMPHOMA, SPLEEN
C2856031|T037|S68.617S|ICD10CM|COMPLETE TRAUMATIC TRANSPHALANGEAL AMPUTATION OF LEFT LITTLE FINGER, SEQUELA|COMPLETE TRAUMATIC TRNSPHAL AMP OF L LITTLE FINGER, SEQUELA
C2873813|T047|D71|ICD10CM|FUNCTIONAL DISORDERS OF POLYMORPHONUCLEAR NEUTROPHILS|CELL MEMBRANE RECEPTOR COMPLEX [CR3] DEFECT
C2873761|T047|D57.01|ICD10CM|HB-SS DISEASE WITH ACUTE CHEST SYNDROME|HB-SS DISEASE WITH ACUTE CHEST SYNDROME
C0238425|T047|D57.00|ICD10CM|HB-SS DISEASE WITH CRISIS, UNSPECIFIED|HB-SS DISEASE WITH CRISIS, UNSPECIFIED
C2873762|T047|D57.02|ICD10CM|HB-SS DISEASE WITH SPLENIC SEQUESTRATION|HB-SS DISEASE WITH SPLENIC SEQUESTRATION
C2886728|T037|T79.2XXA|ICD10CM|TRAUMATIC SECONDARY AND RECURRENT HEMORRHAGE AND SEROMA, INITIAL ENCOUNTER|TRAUMATIC SECONDARY AND RECURRENT HEMOR AND SEROMA, INIT
C2879076|T037|T45.2X2A|ICD10CM|POISONING BY VITAMINS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY VITAMINS, INTENTIONAL SELF-HARM, INIT ENCNTR
C2869761|T037|S98.012S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT FOOT AT ANKLE LEVEL, SEQUELA|COMPLETE TRAUMATIC AMP OF LEFT FOOT AT ANKLE LEVEL, SEQUELA
C0403428|T047|N03.3|DMDICD10|CHRONIC NEPHRITIC SYNDROME WITH DIFFUSE MESANGIAL PROLIFERATIVE GLOMERULONEPHRITIS|CHRONISCHES NEPHRITISCHES SYNDROM: DIFFUSE MESANGIOPROLIFERATIVE GLOMERULONEPHRITIS
C0017665|T047|N03.2|DMDICD10|CHRONIC NEPHRITIC SYNDROME WITH DIFFUSE MEMBRANOUS GLOMERULONEPHRITIS|CHRONISCHES NEPHRITISCHES SYNDROM: DIFFUSE MEMBRANOESE GLOMERULONEPHRITIS
C2902879|T047|N03.1|ICD10CM|CHRONIC NEPHRITIC SYNDROME WITH FOCAL AND SEGMENTAL GLOMERULAR LESIONS|CHRONIC NEPHRITIC SYNDROME WITH FOCAL GLOMERULONEPHRITIS
C2902876|T047|N03.0|ICD10CM|CHRONIC NEPHRITIC SYNDROME WITH MINOR GLOMERULAR ABNORMALITY|CHRONIC NEPHRITIC SYNDROME WITH MINIMAL CHANGE LESION
C2902882|T047|N03.7|ICD10CM|CHRONIC NEPHRITIC SYNDROME WITH DIFFUSE CRESCENTIC GLOMERULONEPHRITIS|CHRONIC NEPHRITIC SYNDROME WITH EXTRACAPILLARY GLOMERULONEPHRITIS
C2902881|T047|N03.6|ICD10CM|CHRONIC NEPHRITIC SYNDROME WITH DENSE DEPOSIT DISEASE|CHRONIC NEPHRITIC SYNDROME WITH MEMBRANOPROLIFERATIVE GLOMERULONEPHRITIS, TYPE 2
C2902880|T047|N03.5|ICD10CM|CHRONIC NEPHRITIC SYNDROME WITH DIFFUSE MESANGIOCAPILLARY GLOMERULONEPHRITIS|CHRONIC NEPHRITIC SYNDROME WITH MEMBRANOPROLIFERATIVE GLOMERULONEPHRITIS, TYPES 1 AND 3, OR NOS
C0451745|T047|N03.4|DMDICD10|CHRONIC NEPHRITIC SYNDROME WITH DIFFUSE ENDOCAPILLARY PROLIFERATIVE GLOMERULONEPHRITIS|CHRONISCHES NEPHRITISCHES SYNDROM: DIFFUSE ENDOKAPILLAER-PROLIFERATIVE GLOMERULONEPHRITIS
C2902885|T047|N03.9|ICD10CM|CHRONIC NEPHRITIC SYNDROME WITH UNSPECIFIED MORPHOLOGIC CHANGES|CHRONIC NEPHRITIC SYNDROME WITH UNSP MORPHOLOGIC CHANGES
C2902884|T047|N03.8|ICD10CM|CHRONIC NEPHRITIC SYNDROME WITH OTHER MORPHOLOGIC CHANGES|CHRONIC NEPHRITIC SYNDROME WITH OTHER MORPHOLOGIC CHANGES
C2890626|T037|T84.122A|ICD10CM|DISPLACEMENT OF INTERNAL FIXATION DEVICE OF BONE OF RIGHT FOREARM, INITIAL ENCOUNTER|DISPLACEMENT OF INT FIX OF BONE OF RIGHT FOREARM, INIT
C2859997|T037|S78.111A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN RIGHT HIP AND KNEE, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMP AT LEVEL BETW R HIP AND KNEE, INIT
C2859998|T037|S78.111D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN RIGHT HIP AND KNEE, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMP AT LEVEL BETW R HIP AND KNEE, SUBS
C4270315|T046|T83.511A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INDWELLING URETHRAL CATHETER, INITIAL ENCOUNTER|I/I REACT D/T INDWELLING URETHRAL CATHETER, INIT
C2832136|T037|S06.320A|ICD10CM|CONTUSION AND LACERATION OF LEFT CEREBRUM WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|CONTUS/LAC LEFT CEREBRUM W/O LOSS OF CONSCIOUSNESS, INIT
C2837677|T037|S32.111B|ICD10CM|MINIMALLY DISPLACED ZONE I FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|MINIMALLY DISPLACED ZONE I FX SACRUM, INIT FOR OPN FX
C2837676|T037|S32.111A|ICD10CM|MINIMALLY DISPLACED ZONE I FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|MINIMALLY DISPLACED ZONE I FRACTURE OF SACRUM, INIT
C2832138|T037|S06.320S|ICD10CM|CONTUSION AND LACERATION OF LEFT CEREBRUM WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|CONTUS/LAC LEFT CEREBRUM W/O LOSS OF CONSCIOUSNESS, SEQUELA
C2890459|T037|T84.031A|ICD10CM|MECHANICAL LOOSENING OF INTERNAL LEFT HIP PROSTHETIC JOINT, INITIAL ENCOUNTER|MECH LOOSENING OF INTERNAL LEFT HIP PROSTHETIC JOINT, INIT
C2833428|T037|S12.351B|ICD10CM|OTHER TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH TRAUM NONDISP SPONDYLOLYSIS OF 4TH CERVCAL VERT, 7THB
C2889004|T047|M02.139|ICD10CM|POSTDYSENTERIC ARTHROPATHY, UNSPECIFIED WRIST|POSTDYSENTERIC ARTHROPATHY, UNSPECIFIED WRIST
C2833427|T037|S12.351A|ICD10CM|OTHER TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH TRAUM NONDISP SPONDYLOLYSIS OF FOURTH CERVCAL VERT, INIT
C2889003|T047|M02.132|ICD10CM|POSTDYSENTERIC ARTHROPATHY, LEFT WRIST|POSTDYSENTERIC ARTHROPATHY, LEFT WRIST
C2889002|T047|M02.131|ICD10CM|POSTDYSENTERIC ARTHROPATHY, RIGHT WRIST|POSTDYSENTERIC ARTHROPATHY, RIGHT WRIST
C2832028|T037|S06.2X4A|ICD10CM|DIFFUSE TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|DIFFUSE TBI W LOC OF 6 HOURS TO 24 HOURS, INIT
C2887818|T047|K51.418|ICD10CM|INFLAMMATORY POLYPS OF COLON WITH OTHER COMPLICATION|INFLAMMATORY POLYPS OF COLON WITH OTHER COMPLICATION
C2887819|T047|K51.419|ICD10CM|INFLAMMATORY POLYPS OF COLON WITH UNSPECIFIED COMPLICATIONS|INFLAMMATORY POLYPS OF COLON WITH UNSPECIFIED COMPLICATIONS
C2887817|T047|K51.414|ICD10CM|INFLAMMATORY POLYPS OF COLON WITH ABSCESS|INFLAMMATORY POLYPS OF COLON WITH ABSCESS
C2887815|T047|K51.412|ICD10CM|INFLAMMATORY POLYPS OF COLON WITH INTESTINAL OBSTRUCTION|INFLAMMATORY POLYPS OF COLON WITH INTESTINAL OBSTRUCTION
C2887816|T047|K51.413|ICD10CM|INFLAMMATORY POLYPS OF COLON WITH FISTULA|INFLAMMATORY POLYPS OF COLON WITH FISTULA
C2887814|T047|K51.411|ICD10CM|INFLAMMATORY POLYPS OF COLON WITH RECTAL BLEEDING|INFLAMMATORY POLYPS OF COLON WITH RECTAL BLEEDING
C2887843|T047|K51.914|ICD10CM|ULCERATIVE COLITIS, UNSPECIFIED WITH ABSCESS|ULCERATIVE COLITIS, UNSPECIFIED WITH ABSCESS
C2832030|T037|S06.2X4S|ICD10CM|DIFFUSE TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|DIFFUSE TBI W LOC OF 6 HOURS TO 24 HOURS, SEQUELA
C0154275|T046|D80.4|DMDICD10|SELECTIVE DEFICIENCY OF IMMUNOGLOBULIN M [IGM]|SELEKTIVER IMMUNGLOBULIN-M-MANGEL [IGM-MANGEL]
C2887841|T047|K51.912|ICD10CM|ULCERATIVE COLITIS, UNSPECIFIED WITH INTESTINAL OBSTRUCTION|ULCERATIVE COLITIS, UNSPECIFIED WITH INTESTINAL OBSTRUCTION
C2832608|T037|S06.824S|ICD10CM|INJURY OF LEFT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|INJURY OF L INT CAROTID, INTCR W LOC OF 6-24 HRS, SEQUELA
C0475535|T047|D80.6|DMDICD10|ANTIBODY DEFICIENCY WITH NEAR-NORMAL IMMUNOGLOBULINS OR WITH HYPERIMMUNOGLOBULINEMIA|ANTIKOERPERMANGEL BEI NORMO- ODER HYPERGAMMAGLOBULINAEMIE
C2882194|T047|I25.750|ICD10CM|ATHEROSCLEROSIS OF NATIVE CORONARY ARTERY OF TRANSPLANTED HEART WITH UNSTABLE ANGINA|ATHSCL NATIVE COR ART OF TXPLT HEART W UNSTABLE ANGINA
C2882195|T047|I25.751|ICD10CM|ATHEROSCLEROSIS OF NATIVE CORONARY ARTERY OF TRANSPLANTED HEART WITH ANGINA PECTORIS WITH DOCUMENTED SPASM|ATHSCL NATIVE COR ART OF TXPLT HEART W ANG PCTRS W SPASM
C0520676|T048||ICD10CM|PREMENSTRUAL DYSPHORIC DISORDER
C2882196|T047|I25.758|ICD10CM|ATHEROSCLEROSIS OF NATIVE CORONARY ARTERY OF TRANSPLANTED HEART WITH OTHER FORMS OF ANGINA PECTORIS|ATHSCL NATIVE COR ART OF TRANSPLANTED HEART W OTH ANG PCTRS
C2882197|T047|I25.759|ICD10CM|ATHEROSCLEROSIS OF NATIVE CORONARY ARTERY OF TRANSPLANTED HEART WITH UNSPECIFIED ANGINA PECTORIS|ATHSCL NATIVE COR ART OF TRANSPLANTED HEART W UNSP ANG PCTRS
C4268302|T048|F32.89|ICD10CM|OTHER SPECIFIED DEPRESSIVE EPISODES|SINGLE EPISODE OF 'MASKED' DEPRESSION NOS
C0348249|T047|B44.89|ICD10CM|OTHER FORMS OF ASPERGILLOSIS|OTHER FORMS OF ASPERGILLOSIS
C0004031|T047||ICD10CM|ALLERGIC BRONCHOPULMONARY ASPERGILLOSIS
C2856982|T037|S72.063A|ICD10CM|DISPLACED ARTICULAR FRACTURE OF HEAD OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED ARTICULAR FRACTURE OF HEAD OF UNSP FEMUR, INIT
C2853718|T191|C81.07|ICD10CM|NODULAR LYMPHOCYTE PREDOMINANT HODGKIN LYMPHOMA, SPLEEN|NODULAR LYMPHOCYTE PREDOMINANT HODGKIN LYMPHOMA, SPLEEN
C2853717|T191|C81.06|ICD10CM|NODULAR LYMPHOCYTE PREDOMINANT HODGKIN LYMPHOMA, INTRAPELVIC LYMPH NODES|NODULAR LYMPHOCYTE PREDOM HODGKIN LYMPHOMA, INTRAPELV NODES
C2853716|T191|C81.05|ICD10CM|NODULAR LYMPHOCYTE PREDOMINANT HODGKIN LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|NODLR LYMPHOCY PREDOM HDGKN LYMPH,NODES OF ING RGN & LOW LMB
C2853715|T191|C81.04|ICD10CM|NODULAR LYMPHOCYTE PREDOMINANT HODGKIN LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB|NODLR LYMPHOCY PREDOM HDGKN LYMPH, NODES OF AXLA AND UPR LMB
C2853714|T191|C81.03|ICD10CM|NODULAR LYMPHOCYTE PREDOMINANT HODGKIN LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES|NODULAR LYMPHOCYTE PREDOM HODGKIN LYMPHOMA, INTRA-ABD NODES
C2853713|T191|C81.02|ICD10CM|NODULAR LYMPHOCYTE PREDOMINANT HODGKIN LYMPHOMA, INTRATHORACIC LYMPH NODES|NODULAR LYMPHOCY PREDOM HODGKIN LYMPHOMA, INTRATHORAC NODES
C2853712|T191|C81.01|ICD10CM|NODULAR LYMPHOCYTE PREDOMINANT HODGKIN LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK|NODLR LYMPHOCY PREDOM HDGKN LYMPH, NODES OF HEAD, FACE, & NK
C2853711|T191|C81.00|ICD10CM|NODULAR LYMPHOCYTE PREDOMINANT HODGKIN LYMPHOMA, UNSPECIFIED SITE|NODULAR LYMPHOCYTE PREDOMINANT HODGKIN LYMPHOMA, UNSP SITE
C2882583|T047|I69.343|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING CEREBRAL INFARCTION AFFECTING RIGHT NON-DOMINANT SIDE|MONOPLG LOW LMB FOL CEREBRAL INFRC AFF RIGHT NONDOM SIDE
C2882582|T047|I69.342|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING CEREBRAL INFARCTION AFFECTING LEFT DOMINANT SIDE|MONOPLG LOW LMB FOL CEREBRAL INFRC AFF LEFT DOMINANT SIDE
C2882581|T047|I69.341|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING CEREBRAL INFARCTION AFFECTING RIGHT DOMINANT SIDE|MONOPLG LOW LMB FOL CEREBRAL INFRC AFF RIGHT DOMINANT SIDE
C2856984|T037|S72.063C|ICD10CM|DISPLACED ARTICULAR FRACTURE OF HEAD OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL ARTIC FX HEAD OF UNSP FEMR, 7THC
C2853720|T191|C81.09|ICD10CM|NODULAR LYMPHOCYTE PREDOMINANT HODGKIN LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES|NODLR LYMPHOCY PREDOM HDGKN LYMPH, EXTRNOD & SOLID ORG SITE
C2853719|T191|C81.08|ICD10CM|NODULAR LYMPHOCYTE PREDOMINANT HODGKIN LYMPHOMA, LYMPH NODES OF MULTIPLE SITES|NODULAR LYMPHOCYTE PREDOM HODGKIN LYMPHOMA, NODES MULT SITE
C2869828|T037|S98.149A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF ONE UNSPECIFIED LESSER TOE, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF ONE UNSP LESSER TOE, INIT
C2889175|T047|M05.231|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT WRIST|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF RIGHT WRIST
C2832407|T037|S06.385A|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF BRAINSTEM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, INITIAL ENCOUNTER|CONTUS/LAC/HEM BRAINSTEM W LOC >24 HR W RET CONSC LEV, INIT
C2888824|T047|M00.079|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, UNSPECIFIED ANKLE AND FOOT|STAPHYLOCOCCAL ARTHRITIS, UNSPECIFIED ANKLE AND FOOT
C2886759|T037|T79.A19A|ICD10CM|TRAUMATIC COMPARTMENT SYNDROME OF UNSPECIFIED UPPER EXTREMITY, INITIAL ENCOUNTER|TRAUMATIC COMPARTMENT SYNDROME OF UNSP UPPER EXTREMITY, INIT
C2888822|T047|M00.071|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, RIGHT ANKLE AND FOOT|STAPHYLOCOCCAL ARTHRITIS, RIGHT ANKLE AND FOOT
C2888823|T047|M00.072|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, LEFT ANKLE AND FOOT|STAPHYLOCOCCAL ARTHRITIS, LEFT ANKLE AND FOOT
C2882809|T047|I70.412|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, LEFT LEG|ATHSCL AUTOL VEIN BYPASS OF EXTRM W INTRMT CLAUD, LEFT LEG
C2832409|T037|S06.385S|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF BRAINSTEM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, SEQUELA|CONTUS/LAC/HEM BRNST W LOC >24 HR W RET CONSC LEV, SEQUELA
C4270246|T046|T83.098A|ICD10CM|OTHER MECHANICAL COMPLICATION OF OTHER URINARY CATHETER, INITIAL ENCOUNTER|MECH COMPL OF OTHER URINARY CATHETER, INITIAL ENCOUNTER
C0477686|T047|M86.8|ICD10CM|OTHER OSTEOMYELITIS, UNSPECIFIED SITES|OTHER OSTEOMYELITIS
C2887098|T047|A41.59|ICD10CM|OTHER GRAM-NEGATIVE SEPSIS|OTHER GRAM-NEGATIVE SEPSIS
C0840005|T047|M86.8X7|ICD10CM|OTHER OSTEOMYELITIS, ANKLE AND FOOT|OTHER OSTEOMYELITIS, ANKLE AND FOOT
C0840004|T047|M86.8X6|ICD10CM|OTHER OSTEOMYELITIS, LOWER LEG|OTHER OSTEOMYELITIS, LOWER LEG
C2901934|T047|M86.8X5|ICD10CM|OTHER OSTEOMYELITIS, THIGH|OTHER OSTEOMYELITIS, THIGH
C0840002|T047|M86.8X4|ICD10CM|OTHER OSTEOMYELITIS, HAND|OTHER OSTEOMYELITIS, HAND
C2887096|T047|A41.52|ICD10CM|SEPSIS DUE TO PSEUDOMONAS|SEPSIS DUE TO PSEUDOMONAS
C2887097|T047|A41.53|ICD10CM|SEPSIS DUE TO SERRATIA|SEPSIS DUE TO SERRATIA
C0036685|T047|A41.50|ICD10CM|GRAM-NEGATIVE SEPSIS, UNSPECIFIED|GRAM-NEGATIVE SEPSIS, UNSPECIFIED
C2887094|T047|A41.51|ICD10CM|SEPSIS DUE TO ESCHERICHIA COLI [E. COLI]|SEPSIS DUE TO ESCHERICHIA COLI [E. COLI]
C2977070|T047|J96.20|ICD10CM|ACUTE AND CHRONIC RESPIRATORY FAILURE, UNSPECIFIED WHETHER WITH HYPOXIA OR HYPERCAPNIA|ACUTE AND CHR RESP FAILURE, UNSP W HYPOXIA OR HYPERCAPNIA
C2977071|T047|J96.21|ICD10CM|ACUTE AND CHRONIC RESPIRATORY FAILURE WITH HYPOXIA|ACUTE AND CHRONIC RESPIRATORY FAILURE WITH HYPOXIA
C2977072|T047|J96.22|ICD10CM|ACUTE AND CHRONIC RESPIRATORY FAILURE WITH HYPERCAPNIA|ACUTE AND CHRONIC RESPIRATORY FAILURE WITH HYPERCAPNIA
C4270565|T046|T85.695A|ICD10CM|OTHER MECHANICAL COMPLICATION OF OTHER NERVOUS SYSTEM DEVICE, IMPLANT OR GRAFT, INITIAL ENCOUNTER|MECH COMPL OF NERVOUS SYS DEVICE, IMPLANT OR GRAFT, INIT
C2833947|T037|S14.128A|ICD10CM|CENTRAL CORD SYNDROME AT C8 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|CENTRAL CORD SYNDROME AT C8, INIT
C2838422|T037|S32.609A|ICD10CM|UNSPECIFIED FRACTURE OF UNSPECIFIED ISCHIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF UNSP ISCHIUM, INIT FOR CLOS FX
C2890929|T037|T85.01XA|ICD10CM|BREAKDOWN (MECHANICAL) OF VENTRICULAR INTRACRANIAL (COMMUNICATING) SHUNT, INITIAL ENCOUNTER|BREAKDOWN OF VENTRICULAR INTRACRANIAL SHUNT, INIT
C2874668|T048|F15.93|ICD10CM|OTHER STIMULANT USE, UNSPECIFIED WITH WITHDRAWAL|OTHER STIMULANT USE, UNSPECIFIED WITH WITHDRAWAL
C4268258|T048|F15.94|ICD10CM|OTHER STIMULANT USE, UNSPECIFIED WITH STIMULANT-INDUCED MOOD DISORDER|AMPHETAMINE OR OTHER STIMULANT-INDUCED BIPOLAR OR RELATED DISORDER, WITHOUT USE DISORDER
C2874678|T048|F15.99|ICD10CM|OTHER STIMULANT USE, UNSPECIFIED WITH UNSPECIFIED STIMULANT-INDUCED DISORDER|OTH STIMULANT USE, UNSP WITH UNSP STIMULANT-INDUCED DISORDER
C2834007|T037|S14.144S|ICD10CM|BROWN-SEQUARD SYNDROME AT C4 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|BROWN-SEQUARD SYNDROME AT C4, SEQUELA
C2874547|T048|F13.282|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED SLEEP DISORDER|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE W SLEEP DISORDER
C2874545|T048|F13.280|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED ANXIETY DISORDER|SEDATV/HYP/ANXIOLYTC DEPENDENCE W ANXIETY DISORDER
C2874546|T048|F13.281|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED SEXUAL DYSFUNCTION|SEDATV/HYP/ANXIOLYTC DEPENDENCE W SEXUAL DYSFUNCTION
C3264460|T047|K75.4|ICD10CM|AUTOIMMUNE HEPATITIS|LUPOID HEPATITIS NEC
C2901806|T047|M86.142|ICD10CM|OTHER ACUTE OSTEOMYELITIS, LEFT HAND|OTHER ACUTE OSTEOMYELITIS, LEFT HAND
C2834005|T037|S14.144A|ICD10CM|BROWN-SEQUARD SYNDROME AT C4 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|BROWN-SEQUARD SYNDROME AT C4, INIT
C4268229|T048|F13.288|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH OTHER SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED DISORDER|SEDATIVE, HYPNOTIC, OR ANXIOLYTIC USE DISORDER, SEVERE, WITH SEDATIVE, HYPNOTIC, OR ANXIOLYTIC-INDUCED MILD NEUROCOGNITIVE DISORDER
C2901805|T047|M86.141|ICD10CM|OTHER ACUTE OSTEOMYELITIS, RIGHT HAND|OTHER ACUTE OSTEOMYELITIS, RIGHT HAND
C2834006|T037|S14.144D|ICD10CM|BROWN-SEQUARD SYNDROME AT C4 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|BROWN-SEQUARD SYNDROME AT C4, SUBS
C2882333|T047|I63.019|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF UNSPECIFIED VERTEBRAL ARTERY|CEREBRAL INFARCTION DUE TO THOMBOS UNSP VERTEBRAL ARTERY
C2890650|T037|T84.129A|ICD10CM|DISPLACEMENT OF INTERNAL FIXATION DEVICE OF UNSPECIFIED BONE OF LIMB, INITIAL ENCOUNTER|DISPLACEMENT OF INT FIX OF UNSP BONE OF LIMB, INIT
C2842081|T191|C50.021|ICD10CM|MALIGNANT NEOPLASM OF NIPPLE AND AREOLA, RIGHT MALE BREAST|MALIGNANT NEOPLASM OF NIPPLE AND AREOLA, RIGHT MALE BREAST
C2889279|T047|M05.541|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT HAND|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT HAND
C2882331|T047|I63.011|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF RIGHT VERTEBRAL ARTERY|CEREBRAL INFARCTION DUE TO THROMBOSIS OF R VERTEB ART
C4268475|T047|I63.013|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF BILATERAL VERTEBRAL ARTERIES|CEREBRAL INFRC DUE TO THROMBOSIS OF BILATERAL VERTEB ART
C2882332|T047|I63.012|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF LEFT VERTEBRAL ARTERY|CEREBRAL INFARCTION DUE TO THROMBOSIS OF L VERTEB ART
C2842083|T191|C50.029|ICD10CM|MALIGNANT NEOPLASM OF NIPPLE AND AREOLA, UNSPECIFIED MALE BREAST|MALIGNANT NEOPLASM OF NIPPLE AND AREOLA, UNSP MALE BREAST
C2889281|T047|M05.549|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP HAND
C3264220|T047|H40.1324|ICD10CM|PIGMENTARY GLAUCOMA, LEFT EYE, INDETERMINATE STAGE|PIGMENTARY GLAUCOMA, LEFT EYE, INDETERMINATE STAGE
C4290152|T047|I70.25|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF OTHER EXTREMITIES WITH ULCERATION|ANY CONDITION CLASSIFIABLE TO I70.218 AND I70.228
C3264217|T047|H40.1321|ICD10CM|PIGMENTARY GLAUCOMA, LEFT EYE, MILD STAGE|PIGMENTARY GLAUCOMA, LEFT EYE, MILD STAGE
C3264216|T047|H40.1320|ICD10CM|PIGMENTARY GLAUCOMA, LEFT EYE, STAGE UNSPECIFIED|PIGMENTARY GLAUCOMA, LEFT EYE, STAGE UNSPECIFIED
C3264219|T047|H40.1323|ICD10CM|PIGMENTARY GLAUCOMA, LEFT EYE, SEVERE STAGE|PIGMENTARY GLAUCOMA, LEFT EYE, SEVERE STAGE
C3264218|T047|H40.1322|ICD10CM|PIGMENTARY GLAUCOMA, LEFT EYE, MODERATE STAGE|PIGMENTARY GLAUCOMA, LEFT EYE, MODERATE STAGE
C2835841|T037|S24.151A|ICD10CM|OTHER INCOMPLETE LESION AT T1 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|OTH INCOMPLETE LESION AT T1, INIT
C2890894|T037|T84.7XXA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO OTHER INTERNAL ORTHOPEDIC PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|INFECT/INFLM REACT DUE TO OTH INT ORTH PROSTH DEV/GRFT, INIT
C0837546|T047|M05.60|ICD10CM|RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF UNSP SITE W INVOLV OF ORGANS AND SYSTEMS
C2833916|T037|S14.119S|ICD10CM|COMPLETE LESION AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, SEQUELA|COMPLETE LESION AT UNSP LEVEL OF CERV SPINAL CORD, SEQUELA
C0837537|T047|M05.69|ICD10CM|RHEUMATOID ARTHRITIS OF MULTIPLE SITES WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS MULT SITE W INVOLV OF ORGANS AND SYSTEMS
C2835843|T037|S24.151S|ICD10CM|OTHER INCOMPLETE LESION AT T1 LEVEL OF THORACIC SPINAL CORD, SEQUELA|OTH INCOMPLETE LESION AT T1, SEQUELA
C2859079|T037|S72.90XA|ICD10CM|UNSPECIFIED FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF UNSP FEMUR, INIT ENCNTR FOR CLOSED FRACTURE
C2859080|T037|S72.90XB|ICD10CM|UNSPECIFIED FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP FRACTURE OF UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2859081|T037|S72.90XC|ICD10CM|UNSPECIFIED FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP FRACTURE OF UNSP FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2833915|T037|S14.119D|ICD10CM|COMPLETE LESION AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION AT UNSP LEVEL OF CERVICAL SPINAL CORD, SUBS
C2833914|T037|S14.119A|ICD10CM|COMPLETE LESION AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION AT UNSP LEVEL OF CERVICAL SPINAL CORD, INIT
C2889333|T047|M05.722|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT ELBOW WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRITIS W RHEU FACTOR OF L ELBOW W/O ORG/SYS INVOLV
C2889332|T047|M05.721|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT ELBOW WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRITIS W RHEU FACTOR OF R ELBOW W/O ORG/SYS INVOLV
C2831613|T037|S02.91XS|ICD10CM|UNSPECIFIED FRACTURE OF SKULL, SEQUELA|UNSPECIFIED FRACTURE OF SKULL, SEQUELA
C4269235|T037|S02.101S|ICD10CM|FRACTURE OF BASE OF SKULL, RIGHT SIDE, SEQUELA|FRACTURE OF BASE OF SKULL, RIGHT SIDE, SEQUELA
C2874376|T048|F10.151|ICD10CM|ALCOHOL ABUSE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|ALCOHOL ABUSE W ALCOH-INDUCE PSYCHOTIC DISORDER W HALLUCIN
C2874375|T048|F10.150|ICD10CM|ALCOHOL ABUSE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|ALCOHOL ABUSE W ALCOH-INDUCE PSYCHOTIC DISORDER W DELUSIONS
C4270196|T046|T83.018A|ICD10CM|BREAKDOWN (MECHANICAL) OF OTHER URINARY CATHETER, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF OTHER URINARY CATHETER, INIT
C4269370|T037|S02.402A|ICD10CM|ZYGOMATIC FRACTURE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|ZYGOMATIC FRACTURE, UNSPECIFIED SIDE, INIT
C2889334|T047|M05.729|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED ELBOW WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRIT W RHEU FACTOR OF UNSP ELBOW W/O ORG/SYS INVOLV
C2874377|T048|F10.159|ICD10CM|ALCOHOL ABUSE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|ALCOHOL ABUSE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED
C2831608|T037|S02.91XA|ICD10CM|UNSPECIFIED FRACTURE OF SKULL, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF SKULL, INIT ENCNTR FOR CLOSED FRACTURE
C2831609|T037|S02.91XB|ICD10CM|UNSPECIFIED FRACTURE OF SKULL, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSPECIFIED FRACTURE OF SKULL, INIT ENCNTR FOR OPEN FRACTURE
C4269231|T037|S02.101B|ICD10CM|FRACTURE OF BASE OF SKULL, RIGHT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF BASE OF SKULL, RIGHT SIDE, 7THB
C2884913|T037|T59.5X2A|ICD10CM|TOXIC EFFECT OF FLUORINE GAS AND HYDROGEN FLUORIDE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOX EFF OF FLUORINE GAS AND HYDROGEN FLUORIDE, SLF-HRM, INIT
C4269230|T037|S02.101A|ICD10CM|FRACTURE OF BASE OF SKULL, RIGHT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF BASE OF SKULL, RIGHT SIDE, INIT
C4269375|T037|S02.402S|ICD10CM|ZYGOMATIC FRACTURE, UNSPECIFIED SIDE, SEQUELA|ZYGOMATIC FRACTURE, UNSPECIFIED SIDE, SEQUELA
C2901567|T046|M84.674A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, RIGHT FOOT, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, RIGHT FOOT, INIT
C2877307|T037|T38.992S|ICD10CM|POISONING BY OTHER HORMONE ANTAGONISTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH HORMONE ANTAGONISTS, SELF-HARM, SEQUELA
C2874947|T048|F40.298|ICD10CM|OTHER SPECIFIED PHOBIA|OTHER SPECIFIED PHOBIA
C2905742|T037|X77.8XXA|ICD10CM|INTENTIONAL SELF-HARM BY OTHER HOT OBJECTS, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY OTHER HOT OBJECTS, INIT ENCNTR
C0522195|T048|F40.291|ICD10CM|GYNEPHOBIA|GYNEPHOBIA
C0522194|T048|F40.290|ICD10CM|ANDROPHOBIA|ANDROPHOBIA
C2890357|T037|T83.498A|ICD10CM|OTHER MECHANICAL COMPLICATION OF OTHER PROSTHETIC DEVICES, IMPLANTS AND GRAFTS OF GENITAL TRACT, INITIAL ENCOUNTER|MECH COMPL OF PROSTH DEV/IMPLNT/GRFT OF GENITAL TRACT, INIT
C2877305|T037|T38.992A|ICD10CM|POISONING BY OTHER HORMONE ANTAGONISTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH HORMONE ANTAGONISTS, SELF-HARM, INIT
C2012187|T047||ICD10CM|RESIDUAL STAGE OF OPEN-ANGLE GLAUCOMA, RIGHT EYE
C2012186|T047||ICD10CM|RESIDUAL STAGE OF OPEN-ANGLE GLAUCOMA, LEFT EYE
C2881011|T047|H40.153|ICD10CM|RESIDUAL STAGE OF OPEN-ANGLE GLAUCOMA, BILATERAL|RESIDUAL STAGE OF OPEN-ANGLE GLAUCOMA, BILATERAL
C2900947|T046|M84.441A|ICD10CM|PATHOLOGICAL FRACTURE, RIGHT HAND, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, RIGHT HAND, INIT ENCNTR FOR FRACTURE
C2881012|T047|H40.159|ICD10CM|RESIDUAL STAGE OF OPEN-ANGLE GLAUCOMA, UNSPECIFIED EYE|RESIDUAL STAGE OF OPEN-ANGLE GLAUCOMA, UNSPECIFIED EYE
C2890247|T037|T83.111A|ICD10CM|BREAKDOWN (MECHANICAL) OF IMPLANTED URINARY SPHINCTER, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF IMPLANTED URINARY SPHINCTER, INIT
C2860064|T037|S79.009A|ICD10CM|UNSPECIFIED PHYSEAL FRACTURE OF UPPER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP PHYSEAL FRACTURE OF UPPER END OF UNSP FEMUR, INIT
C2887480|T046|J68.4|ICD10CM|CHRONIC RESPIRATORY CONDITIONS DUE TO CHEMICALS, GASES, FUMES AND VAPORS|PULMONARY FIBROSIS (CHRONIC) DUE TO INHALATION OF CHEMICALS, GASES, FUMES AND VAPORS
C0494670|T047|J68.0|DMDICD10|BRONCHITIS AND PNEUMONITIS DUE TO CHEMICALS, GASES, FUMES AND VAPORS|BRONCHITIS UND PNEUMONIE DURCH CHEMISCHE SUBSTANZEN, GASE, RAUCH UND DAEMPFE
C2887477|T047|J68.1|ICD10CM|PULMONARY EDEMA DUE TO CHEMICALS, GASES, FUMES AND VAPORS|PULMONARY EDEMA DUE TO CHEMICALS, GASES, FUMES AND VAPORS
C1144817|T047|J68.2|ICD10CM|UPPER RESPIRATORY INFLAMMATION DUE TO CHEMICALS, GASES, FUMES AND VAPORS, NOT ELSEWHERE CLASSIFIED|UPPER RESP INFLAM D/T CHEMICALS, GAS, FUMES AND VAPORS, NEC
C1299633|T047|J68.3|ICD10CM|OTHER ACUTE AND SUBACUTE RESPIRATORY CONDITIONS DUE TO CHEMICALS, GASES, FUMES AND VAPORS|REACTIVE AIRWAYS DYSFUNCTION SYNDROME
C4268014|T047|E10.3219|ICD10CM|TYPE 1 DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|TYPE 1 DIAB WITH MILD NONP RTNOP WITH MACULAR EDEMA, UNSP
C0348700|T046|J68.8|DMDICD10|OTHER RESPIRATORY CONDITIONS DUE TO CHEMICALS, GASES, FUMES AND VAPORS|SONSTIGE KRANKHEITEN DER ATMUNGSORGANE DURCH CHEMISCHE SUBSTANZEN, GASE, RAUCH UND DAEMPFE
C0494673|T047|J68.9|DMDICD10|UNSPECIFIED RESPIRATORY CONDITION DUE TO CHEMICALS, GASES, FUMES AND VAPORS|NICHT NAEHER BEZEICHNETE KRANKHEIT DER ATMUNGSORGANE DURCH CHEMISCHE SUBSTANZEN, GASE, RAUCH UND DAEMPFE
C2902114|T046|M87.365|ICD10CM|OTHER SECONDARY OSTEONECROSIS, LEFT FIBULA|OTHER SECONDARY OSTEONECROSIS, LEFT FIBULA
C2842124|T191|C50.622|ICD10CM|MALIGNANT NEOPLASM OF AXILLARY TAIL OF LEFT MALE BREAST|MALIGNANT NEOPLASM OF AXILLARY TAIL OF LEFT MALE BREAST
C2902115|T046|M87.366|ICD10CM|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED FIBULA|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED FIBULA
C2902110|T046|M87.361|ICD10CM|OTHER SECONDARY OSTEONECROSIS, RIGHT TIBIA|OTHER SECONDARY OSTEONECROSIS, RIGHT TIBIA
C2902112|T046|M87.363|ICD10CM|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED TIBIA|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED TIBIA
C2902111|T046|M87.362|ICD10CM|OTHER SECONDARY OSTEONECROSIS, LEFT TIBIA|OTHER SECONDARY OSTEONECROSIS, LEFT TIBIA
C1318550|T191||ICD10CM|REFRACTORY ANEMIA WITH EXCESS OF BLASTS 1
C0002894|T191|D46.20|ICD10CM|REFRACTORY ANEMIA WITH EXCESS OF BLASTS, UNSPECIFIED|REFRACTORY ANEMIA WITH EXCESS OF BLASTS, UNSPECIFIED
C1318551|T191||ICD10CM|REFRACTORY ANEMIA WITH EXCESS OF BLASTS 2
C4268048|T047|E10.3539|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, UNSPECIFIED EYE|TYPE 1 DIAB W PROLIF DIAB RTNOP WITH TRCTN DTCH N-MCLA, UNSP
C2890336|T037|T83.418A|ICD10CM|BREAKDOWN (MECHANICAL) OF OTHER PROSTHETIC DEVICES, IMPLANTS AND GRAFTS OF GENITAL TRACT, INITIAL ENCOUNTER|BREAKDOWN OF PROSTH DEV/IMPLNT/GRFT OF GENITL TRCT, INIT
C4268045|T047|E10.3531|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, RIGHT EYE|TYPE 1 DIAB W PROLIF DIAB RTNOP W TRCTN DTCH N-MCLA, R EYE
C4268046|T047|E10.3532|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, LEFT EYE|TYPE 1 DIAB W PROLIF DIAB RTNOP W TRCTN DTCH N-MCLA, L EYE
C4268047|T047|E10.3533|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, BILATERAL|TYPE 1 DIAB W PROLIF DIAB RTNOP WITH TRCTN DTCH N-MCLA, BI
C4270173|T046|T82.858A|ICD10CM|STENOSIS OF OTHER VASCULAR PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|STENOSIS OF OTHER VASCULAR PROSTH DEV/GRFT, INIT
C4268011|T047|E10.3211|ICD10CM|TYPE 1 DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|TYPE 1 DIAB WITH MILD NONP RTNOP WITH MACULAR EDEMA, R EYE
C2838700|T037|S34.132S|ICD10CM|INCOMPLETE LESION OF SACRAL SPINAL CORD, SEQUELA|INCOMPLETE LESION OF SACRAL SPINAL CORD, SEQUELA
C2858629|T037|S72.436C|ICD10CM|NONDISPLACED FRACTURE OF MEDIAL CONDYLE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF MED CONDYLE OF UNSP FEMR, 7THC
C2858627|T037|S72.436A|ICD10CM|NONDISPLACED FRACTURE OF MEDIAL CONDYLE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF MEDIAL CONDYLE OF UNSP FEMUR, INIT FOR CLOS FX
C4269287|T037|S02.11BB|ICD10CM|TYPE I OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE I OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, 7THB
C2874449|T048|F11.281|ICD10CM|OPIOID DEPENDENCE WITH OPIOID-INDUCED SEXUAL DYSFUNCTION|OPIOID DEPENDENCE WITH OPIOID-INDUCED SEXUAL DYSFUNCTION
C2874450|T048|F11.282|ICD10CM|OPIOID DEPENDENCE WITH OPIOID-INDUCED SLEEP DISORDER|OPIOID DEPENDENCE WITH OPIOID-INDUCED SLEEP DISORDER
C2838699|T037|S34.132D|ICD10CM|INCOMPLETE LESION OF SACRAL SPINAL CORD, SUBSEQUENT ENCOUNTER|INCOMPLETE LESION OF SACRAL SPINAL CORD, SUBS ENCNTR
C2874448|T048|F11.288|ICD10CM|OPIOID DEPENDENCE WITH OTHER OPIOID-INDUCED DISORDER|OPIOID DEPENDENCE WITH OTHER OPIOID-INDUCED DISORDER
C2885493|T037|T63.192S|ICD10CM|TOXIC EFFECT OF VENOM OF OTHER REPTILES, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF REPTILES, SELF-HARM, SEQUELA
C2838698|T037|S34.132A|ICD10CM|INCOMPLETE LESION OF SACRAL SPINAL CORD, INITIAL ENCOUNTER|INCOMPLETE LESION OF SACRAL SPINAL CORD, INITIAL ENCOUNTER
C2878921|T037|T44.7X2A|ICD10CM|POISONING BY BETA-ADRENORECEPTOR ANTAGONISTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY BETA-ADRENOCPT ANTAGONISTS, SELF-HARM, INIT
C2885731|T037|T63.512S|ICD10CM|TOXIC EFFECT OF CONTACT WITH STINGRAY, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CONTACT W STINGRAY, SELF-HARM, SEQUELA
C2842125|T191|C50.629|ICD10CM|MALIGNANT NEOPLASM OF AXILLARY TAIL OF UNSPECIFIED MALE BREAST|MALIGNANT NEOPLASM OF AXILLARY TAIL OF UNSP MALE BREAST
C2869893|T037|S98.912S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT FOOT, LEVEL UNSPECIFIED, SEQUELA|COMPLETE TRAUMATIC AMP OF LEFT FOOT, LEVEL UNSP, SEQUELA
C0477676|T047|M83.8|DMDICD10|OTHER ADULT OSTEOMALACIA|SONSTIGE OSTEOMALAZIE IM ERWACHSENENALTER
C2883019|T047|I70.763|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, BILATERAL LEGS|ATHSCL TYPE OF BYPASS OF THE EXTRM W GANGRENE, BI LEGS
C2883018|T047|I70.762|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, LEFT LEG|ATHSCL TYPE OF BYPASS OF THE EXTRM W GANGRENE, LEFT LEG
C2883017|T047|I70.761|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, RIGHT LEG|ATHSCL TYPE OF BYPASS OF THE EXTRM W GANGRENE, RIGHT LEG
C2885729|T037|T63.512A|ICD10CM|TOXIC EFFECT OF CONTACT WITH STINGRAY, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CONTACT W STINGRAY, SELF-HARM, INIT
C2874702|T048|F16.259|ICD10CM|HALLUCINOGEN DEPENDENCE WITH HALLUCINOGEN-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|HALLUCINOGEN DEPENDENCE WITH HALLUCINOGEN-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED
C2837730|T037|S32.130B|ICD10CM|NONDISPLACED ZONE III FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISPLACED ZONE III FRACTURE OF SACRUM, INIT FOR OPN FX
C2883021|T047|I70.769|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, UNSPECIFIED EXTREMITY|ATHSCL TYPE OF BYPASS OF THE EXTRM W GANGRENE, UNSP EXTRM
C2883020|T047|I70.768|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, OTHER EXTREMITY|ATHSCL TYPE OF BYPASS OF THE EXTRM W GANGRENE, OTH EXTREMITY
C2874700|T048|F16.250|ICD10CM|HALLUCINOGEN DEPENDENCE WITH HALLUCINOGEN-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|HALLUCINOGEN DEPENDENCE W PSYCHOTIC DISORDER W DELUSIONS
C2874701|T048|F16.251|ICD10CM|HALLUCINOGEN DEPENDENCE WITH HALLUCINOGEN-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|HALLUCINOGEN DEPENDENCE W PSYCHOTIC DISORDER W HALLUCIN
C2884302|T037|T53.6X2A|ICD10CM|TOXIC EFFECT OF OTHER HALOGEN DERIVATIVES OF ALIPHATIC HYDROCARBONS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOX EFF OF HALGN DERIV OF ALIPHATIC HYDROCRB, SLF-HRM, INIT
C0477680|T047|M83|DMDICD10|ADULT OSTEOMALACIA, UNSPECIFIED|OSTEOMALAZIE IM ERWACHSENENALTER
C0153678|T191|C78.2|DMDICD10|SECONDARY MALIGNANT NEOPLASM OF PLEURA|SEKUNDAERE BOESARTIGE NEUBILDUNG DER PLEURA
C0153677|T191|C78.1|DMDICD10|SECONDARY MALIGNANT NEOPLASM OF MEDIASTINUM|SEKUNDAERE BOESARTIGE NEUBILDUNG DES MEDIASTINUMS
C0036528|T191|C78.6|DMDICD10|SECONDARY MALIGNANT NEOPLASM OF RETROPERITONEUM AND PERITONEUM|SEKUNDAERE BOESARTIGE NEUBILDUNG DES RETROPERITONEUMS UND DES PERITONEUMS
C0153364|T191|C03.9|DMDICD10|MALIGNANT NEOPLASM OF GUM, UNSPECIFIED|BOESARTIGE NEUBILDUNG: ZAHNFLEISCH, NICHT NAEHER BEZEICHNET
C0494164|T191|C78.4|DMDICD10|SECONDARY MALIGNANT NEOPLASM OF SMALL INTESTINE|SEKUNDAERE BOESARTIGE NEUBILDUNG DES DUENNDARMES
C0153681|T191|C78.5|DMDICD10|SECONDARY MALIGNANT NEOPLASM OF LARGE INTESTINE AND RECTUM|SEKUNDAERE BOESARTIGE NEUBILDUNG DES DICKDARMES UND DES REKTUMS
C2884304|T037|T53.6X2S|ICD10CM|TOXIC EFFECT OF OTHER HALOGEN DERIVATIVES OF ALIPHATIC HYDROCARBONS, INTENTIONAL SELF-HARM, SEQUELA|TOX EFF OF HALGN DERIV OF ALIPHATIC HYDROCRB, SLF-HRM, SQLA
C2889011|T047|M02.152|ICD10CM|POSTDYSENTERIC ARTHROPATHY, LEFT HIP|POSTDYSENTERIC ARTHROPATHY, LEFT HIP
C2521553|T060|C030|ICD10PCS|MALIGNANT NEOPLASM OF UPPER GUM|NUCLEAR MEDICINE @ CENTRAL NERVOUS SYSTEM @ POSITRON EMISSION TOMOGRAPHIC (PET) IMAGING @ BRAIN
C0432581|T191|C03.1|DMDICD10|MALIGNANT NEOPLASM OF LOWER GUM|BOESARTIGE NEUBILDUNG: UNTERKIEFERZAHNFLEISCH
C2854058|T191|C85.94|ICD10CM|NON-HODGKIN LYMPHOMA, UNSPECIFIED, LYMPH NODES OF AXILLA AND UPPER LIMB|NON-HODGKIN LYMPHOMA, UNSP, NODES OF AXILLA AND UPPER LIMB
C2854059|T191|C85.95|ICD10CM|NON-HODGKIN LYMPHOMA, UNSPECIFIED, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|NON-HODG LYMPHOMA, UNSP, NODES OF ING REGION AND LOWER LIMB
C2854060|T191|C85.96|ICD10CM|NON-HODGKIN LYMPHOMA, UNSPECIFIED, INTRAPELVIC LYMPH NODES|NON-HODGKIN LYMPHOMA, UNSPECIFIED, INTRAPELVIC LYMPH NODES
C2854061|T191|C85.97|ICD10CM|NON-HODGKIN LYMPHOMA, UNSPECIFIED, SPLEEN|NON-HODGKIN LYMPHOMA, UNSPECIFIED, SPLEEN
C2854054|T191|C85.90|ICD10CM|NON-HODGKIN LYMPHOMA, UNSPECIFIED, UNSPECIFIED SITE|NON-HODGKIN LYMPHOMA, UNSPECIFIED, UNSPECIFIED SITE
C4267920|T047|E08.3499|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|DIABETES WITH SEVERE NONP RTNOP WITHOUT MACULAR EDEMA, UNSP
C2854056|T191|C85.92|ICD10CM|NON-HODGKIN LYMPHOMA, UNSPECIFIED, INTRATHORACIC LYMPH NODES|NON-HODGKIN LYMPHOMA, UNSPECIFIED, INTRATHORACIC LYMPH NODES
C2854057|T191|C85.93|ICD10CM|NON-HODGKIN LYMPHOMA, UNSPECIFIED, INTRA-ABDOMINAL LYMPH NODES|NON-HODGKIN LYMPHOMA, UNSP, INTRA-ABDOMINAL LYMPH NODES
C2857841|T037|S72.332C|ICD10CM|DISPLACED OBLIQUE FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL OBLIQUE FX SHAFT OF L FEMR, 7THC
C2857840|T037|S72.332B|ICD10CM|DISPLACED OBLIQUE FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL OBLIQUE FX SHAFT OF L FEMUR, INIT FOR OPN FX TYPE I/2
C2857839|T037|S72.332A|ICD10CM|DISPLACED OBLIQUE FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED OBLIQUE FRACTURE OF SHAFT OF LEFT FEMUR, INIT
C2854062|T191|C85.98|ICD10CM|NON-HODGKIN LYMPHOMA, UNSPECIFIED, LYMPH NODES OF MULTIPLE SITES|NON-HODGKIN LYMPHOMA, UNSP, LYMPH NODES OF MULTIPLE SITES
C2854063|T191|C85.99|ICD10CM|NON-HODGKIN LYMPHOMA, UNSPECIFIED, EXTRANODAL AND SOLID ORGAN SITES|NON-HODGKIN LYMPHOMA, UNSP, EXTRANODAL AND SOLID ORGAN SITES
C4267918|T047|E08.3492|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|DIAB WITH SEVERE NONP RTNOP WITHOUT MACULAR EDEMA, LEFT EYE
C4267919|T047|E08.3493|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|DIABETES WITH SEVERE NONP RTNOP WITHOUT MACULAR EDEMA, BI
C0349053|T191|C25.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF PANCREAS|BOESARTIGE NEUBILDUNG: PANKREAS, MEHRERE TEILBEREICHE UEBERLAPPEND
C0346647|T191|C25.9|DMDICD10|MALIGNANT NEOPLASM OF PANCREAS, UNSPECIFIED|BOESARTIGE NEUBILDUNG: PANKREAS, NICHT NAEHER BEZEICHNET
C0153458|T191|C25.0|DMDICD10|MALIGNANT NEOPLASM OF HEAD OF PANCREAS|BOESARTIGE NEUBILDUNG: PANKREASKOPF
C0153459|T191|C25.1|DMDICD10|MALIGNANT NEOPLASM OF BODY OF PANCREAS|BOESARTIGE NEUBILDUNG: PANKREASKOERPER
C0153460|T191|C25.2|DMDICD10|MALIGNANT NEOPLASM OF TAIL OF PANCREAS|BOESARTIGE NEUBILDUNG: PANKREASSCHWANZ
C0153461|T191|C25.3|DMDICD10|MALIGNANT NEOPLASM OF PANCREATIC DUCT|BOESARTIGE NEUBILDUNG: DUCTUS PANCREATICUS
C1328479|T191||ICD10CM|MALIGNANT NEOPLASM OF ENDOCRINE PANCREAS
C2837940|T191|C25.7|ICD10CM|MALIGNANT NEOPLASM OF OTHER PARTS OF PANCREAS|MALIGNANT NEOPLASM OF NECK OF PANCREAS
C2838028|T037|S32.414A|ICD10CM|NONDISPLACED FRACTURE OF ANTERIOR WALL OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF ANTERIOR WALL OF RIGHT ACETABULUM, INIT
C2876569|T037|T36.1X2A|ICD10CM|POISONING BY CEPHALOSPORINS AND OTHER BETA-LACTAM ANTIBIOTICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY CEPHALOSPOR/OTH BETA-LACTM ANTIBIOT, SLF-HRM, INIT
C2832491|T037|S06.5X5S|ICD10CM|TRAUMATIC SUBDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, SEQUELA|TRAUM SUBDR HEM W LOC >24 HR W RET CONSC LEV, SEQUELA
C2838379|T037|S32.511A|ICD10CM|FRACTURE OF SUPERIOR RIM OF RIGHT PUBIS, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF SUPERIOR RIM OF RIGHT PUBIS, INIT FOR CLOS FX
C2876571|T037|T36.1X2S|ICD10CM|POISONING BY CEPHALOSPORINS AND OTHER BETA-LACTAM ANTIBIOTICS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY CEPHALOSPOR/OTH BETA-LACTM ANTIBIOT, SLF-HRM, SQLA
C2832489|T037|S06.5X5A|ICD10CM|TRAUMATIC SUBDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, INITIAL ENCOUNTER|TRAUM SUBDR HEM W LOC >24 HR W RET CONSC LEV, INIT
C2895173|T047|M32.14|ICD10CM|GLOMERULAR DISEASE IN SYSTEMIC LUPUS ERYTHEMATOSUS|GLOMERULAR DISEASE IN SYSTEMIC LUPUS ERYTHEMATOSUS
C2895174|T047|M32.15|ICD10CM|TUBULO-INTERSTITIAL NEPHROPATHY IN SYSTEMIC LUPUS ERYTHEMATOSUS|TUBULO-INTERSTITIAL NEUROPATH IN SYS LUPUS ERYTHEMATOSUS
C2895168|T047|M32.10|ICD10CM|SYSTEMIC LUPUS ERYTHEMATOSUS, ORGAN OR SYSTEM INVOLVEMENT UNSPECIFIED|SYSTEMIC LUPUS ERYTHEMATOSUS, ORGAN OR SYSTEM INVOLV UNSP
C2895169|T047|M32.11|ICD10CM|ENDOCARDITIS IN SYSTEMIC LUPUS ERYTHEMATOSUS|ENDOCARDITIS IN SYSTEMIC LUPUS ERYTHEMATOSUS
C1141942|T047||ICD10CM|PERICARDITIS IN SYSTEMIC LUPUS ERYTHEMATOSUS
C2895171|T047||ICD10CM|LUNG INVOLVEMENT IN SYSTEMIC LUPUS ERYTHEMATOSUS
C2832244|T037|S06.346A|ICD10CM|TRAUMATIC HEMORRHAGE OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|TRAUM HEMOR R CEREB W LOC >24 HR W/O RET CONSC W SURV, INIT
C2895175|T047|M32.19|ICD10CM|OTHER ORGAN OR SYSTEM INVOLVEMENT IN SYSTEMIC LUPUS ERYTHEMATOSUS|OTH ORGAN OR SYSTEM INVOLV IN SYSTEMIC LUPUS ERYTHEMATOSUS
C2888246|T047|L89.023|ICD10CM|PRESSURE ULCER OF LEFT ELBOW, STAGE 3|PRESSURE ULCER OF LEFT ELBOW, STAGE 3
C2888243|T047|L89.022|ICD10CM|PRESSURE ULCER OF LEFT ELBOW, STAGE 2|PRESSURE ULCER OF LEFT ELBOW, STAGE 2
C2888240|T047|L89.021|ICD10CM|PRESSURE ULCER OF LEFT ELBOW, STAGE 1|PRESSURE ULCER OF LEFT ELBOW, STAGE 1
C2888237|T047||ICD10CM|PRESSURE ULCER OF LEFT ELBOW, UNSTAGEABLE
C2865517|T037|S88.011D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT KNEE LEVEL, RIGHT LOWER LEG, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION AT KNEE LEVEL, R LOW LEG, SUBS
C2888249|T047|L89.024|ICD10CM|PRESSURE ULCER OF LEFT ELBOW, STAGE 4|PRESSURE ULCER OF LEFT ELBOW, STAGE 4
C4509274|T047|L89.029|ICD10CM|PRESSURE ULCER OF LEFT ELBOW, UNSPECIFIED STAGE|HEALING PRESSURE ULCER OF LEFT ELBOW, UNSPECIFIED STAGE
C2832246|T037|S06.346S|ICD10CM|TRAUMATIC HEMORRHAGE OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|TRAUM HEMOR R CEREB W LOC >24 HR W/O RET CONSC W SURV, SQLA
C2873951|T047|E09.01|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH HYPEROSMOLARITY WITH COMA|DRUG/CHEM DIABETES MELLITUS W HYPEROSMOLARITY W COMA
C2873950|T047|E09.00|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH HYPEROSMOLARITY WITHOUT NONKETOTIC HYPERGLYCEMIC-HYPEROSMOLAR COMA (NKHHC)|DRUG/CHEM DIAB W HYPROSM W/O NONKET HYPRGLY-HYPROS COMA
C2889475|T047|M06.831|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, RIGHT WRIST|OTHER SPECIFIED RHEUMATOID ARTHRITIS, RIGHT WRIST
C2885628|T037|T63.422S|ICD10CM|TOXIC EFFECT OF VENOM OF ANTS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF ANTS, SELF-HARM, SEQUELA
C4269483|T037|S02.630B|ICD10CM|FRACTURE OF CORONOID PROCESS OF MANDIBLE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FX CORONOID PROCESS OF MANDIBLE, UNSPECIFIED SIDE, 7THB
C4269482|T037|S02.630A|ICD10CM|FRACTURE OF CORONOID PROCESS OF MANDIBLE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FX CORONOID PROCESS OF MANDIBLE, UNSPECIFIED SIDE, INIT
C2856862|T037|S72.045B|ICD10CM|NONDISPLACED FRACTURE OF BASE OF NECK OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF BASE OF NK OF L FEMR, INIT FOR OPN FX TYPE I/2
C2857770|T037|S72.324A|ICD10CM|NONDISPLACED TRANSVERSE FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP TRANSVERSE FRACTURE OF SHAFT OF RIGHT FEMUR, INIT
C2883456|T037|T49.7X2A|ICD10CM|POISONING BY DENTAL DRUGS, TOPICALLY APPLIED, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY DENTAL DRUGS, TOPICALLY APPLIED, SELF-HARM, INIT
C2856863|T037|S72.045C|ICD10CM|NONDISPLACED FRACTURE OF BASE OF NECK OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF BASE OF NK OF L FEMR, 7THC
C4269487|T037|S02.630S|ICD10CM|FRACTURE OF CORONOID PROCESS OF MANDIBLE, UNSPECIFIED SIDE, SEQUELA|FX CORONOID PROCESS OF MANDIBLE, UNSPECIFIED SIDE, SEQUELA
C2901878|T047|M86.442|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, LEFT HAND|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, LEFT HAND
C2901877|T047|M86.441|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, RIGHT HAND|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, RIGHT HAND
C2838064|T037|S32.423A|ICD10CM|DISPLACED FRACTURE OF POSTERIOR WALL OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF POSTERIOR WALL OF UNSP ACETABULUM, INIT
C2838065|T037|S32.423B|ICD10CM|DISPLACED FRACTURE OF POSTERIOR WALL OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISP FX OF POSTERIOR WALL OF UNSP ACETAB, INIT FOR OPN FX
C2901879|T047|M86.449|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, UNSPECIFIED HAND|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, UNSPECIFIED HAND
C0153567|T191|C55|DMDICD10|MALIGNANT NEOPLASM OF UTERUS, PART UNSPECIFIED|BOESARTIGE NEUBILDUNG DES UTERUS, TEIL NICHT NAEHER BEZEICHNET
C0042237|T191|C52|DMDICD10|MALIGNANT NEOPLASM OF VAGINA|BOESARTIGE NEUBILDUNG DER VAGINA
C0153572|T191|C58|DMDICD10|MALIGNANT NEOPLASM OF PLACENTA|BOESARTIGE NEUBILDUNG DER PLAZENTA
C2874451|T048|F11.29|ICD10CM|OPIOID DEPENDENCE WITH UNSPECIFIED OPIOID-INDUCED DISORDER|OPIOID DEPENDENCE WITH UNSPECIFIED OPIOID-INDUCED DISORDER
C2835384|T037|S22.062A|ICD10CM|UNSTABLE BURST FRACTURE OF T7-T8 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSTABLE BURST FRACTURE OF T7-T8 VERTEBRA, INIT FOR CLOS FX
C2874442|T048|F11.23|ICD10CM|OPIOID DEPENDENCE WITH WITHDRAWAL|OPIOID DEPENDENCE WITH WITHDRAWAL
C2882754|T047|I70.313|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, BILATERAL LEGS|ATHSCL UNSP TYPE BYPASS OF THE EXTRM W INTRMT CLAUD, BI LEGS
C4509043|T048|F11.21|ICD10CM|OPIOID DEPENDENCE, IN REMISSION|OPIOID USE DISORDER, SEVERE, IN SUSTAINED REMISSION
C4237239|T048|F11.20|ICD10CM|OPIOID DEPENDENCE, UNCOMPLICATED|OPIOID USE DISORDER, SEVERE
C2835385|T037|S22.062B|ICD10CM|UNSTABLE BURST FRACTURE OF T7-T8 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSTABLE BURST FRACTURE OF T7-T8 VERTEBRA, INIT FOR OPN FX
C4268216|T048|F11.24|ICD10CM|OPIOID DEPENDENCE WITH OPIOID-INDUCED MOOD DISORDER|OPIOID USE DISORDER, MODERATE, WITH OPIOID INDUCED DEPRESSIVE DISORDER
C4269378|T037|S02.40AB|ICD10CM|MALAR FRACTURE, RIGHT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|MALAR FRACTURE, RIGHT SIDE, 7THB
C2860230|T037|S79.191A|ICD10CM|OTHER PHYSEAL FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH PHYSEAL FRACTURE OF LOWER END OF RIGHT FEMUR, INIT
C2901917|T047|M86.622|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, LEFT  HUMERUS|OTHER CHRONIC OSTEOMYELITIS, LEFT HUMERUS
C2888859|T047|M00.20|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, UNSPECIFIED JOINT|OTHER STREPTOCOCCAL ARTHRITIS, UNSPECIFIED JOINT
C2874602|T048|F14.280|ICD10CM|COCAINE DEPENDENCE WITH COCAINE-INDUCED ANXIETY DISORDER|COCAINE DEPENDENCE WITH COCAINE-INDUCED ANXIETY DISORDER
C2267227|T048|F50.2|DMDICD10|BULIMIA NERVOSA|BULIMIA NERVOSA
C2888891|T047|M00.28|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, VERTEBRAE|OTHER STREPTOCOCCAL ARTHRITIS, VERTEBRAE
C2888892|T047|M00.29|ICD10CM|OTHER STREPTOCOCCAL POLYARTHRITIS|OTHER STREPTOCOCCAL POLYARTHRITIS
C1395047|T047||ICD10CM|MYOCARDIAL DEGENERATION
C0264852|T047||ICD10CM|MYOCARDITIS, UNSPECIFIED
C0494599|T046|I51.1|DMDICD10|RUPTURE OF CHORDAE TENDINEAE, NOT ELSEWHERE CLASSIFIED|RUPTUR DER CHORDAE TENDINEAE, ANDERENORTS NICHT KLASSIFIZIERT
C0494600|T020|I51.2|DMDICD10|RUPTURE OF PAPILLARY MUSCLE, NOT ELSEWHERE CLASSIFIED|PAPILLARMUSKELRUPTUR, ANDERENORTS NICHT KLASSIFIZIERT
C0024117|T047|J44.9|DMDICD10|CHRONIC OBSTRUCTIVE PULMONARY DISEASE, UNSPECIFIED|CHRONISCHE OBSTRUKTIVE LUNGENKRANKHEIT, NICHT NAEHER BEZEICHNET
C2889566|T047|M08.26|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, UNSPECIFIED KNEE|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, KNEE
C0348802|T047|B46.1|DMDICD10|RHINOCEREBRAL MUCORMYCOSIS|RHINOZEREBRALE MUKORMYKOSE
C2889567|T047|M08.261|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, RIGHT KNEE|JUVENILE RHEUMATOID ARTHRITIS W SYSTEMIC ONSET, RIGHT KNEE
C2889568|T047|M08.262|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, LEFT KNEE|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, LEFT KNEE
C4268181|T047|E13.37X9|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, UNSPECIFIED EYE|OTH DIAB WITH DIAB MACULAR EDEMA, RESOLVED FOL TRTMT, UNSP
C2879973|T037|T48.202A|ICD10CM|POISONING BY UNSPECIFIED DRUGS ACTING ON MUSCLES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY UNSP DRUGS ACTING ON MUSCLES, SELF-HARM, INIT
C2888877|T047|M00.249|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, UNSPECIFIED HAND|OTHER STREPTOCOCCAL ARTHRITIS, UNSPECIFIED HAND
C2857257|T037|S72.121A|ICD10CM|DISPLACED FRACTURE OF LESSER TROCHANTER OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF LESSER TROCHANTER OF RIGHT FEMUR, INIT
C4268178|T047|E13.37X1|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, RIGHT EYE|OTH DIAB WITH DIAB MACULAR EDEMA, RESOLVED FOL TRTMT, R EYE
C4268179|T047|E13.37X2|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, LEFT EYE|OTH DIAB WITH DIAB MACULAR EDEMA, RESOLVED FOL TRTMT, L EYE
C4268180|T047|E13.37X3|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, BILATERAL|OTH DIAB WITH DIABETIC MACULAR EDEMA, RESOLVED FOL TRTMT, BI
C2888876|T047|M00.242|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, LEFT HAND|OTHER STREPTOCOCCAL ARTHRITIS, LEFT HAND
C2888875|T047|M00.241|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, RIGHT HAND|OTHER STREPTOCOCCAL ARTHRITIS, RIGHT HAND
C2887468|T047|J47.0|ICD10CM|BRONCHIECTASIS WITH ACUTE LOWER RESPIRATORY INFECTION|BRONCHIECTASIS WITH ACUTE LOWER RESPIRATORY INFECTION
C2882304|T047|I60.32|ICD10CM|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM LEFT POSTERIOR COMMUNICATING ARTERY|NTRM SUBARACH HEMOR FROM LEFT POSTERIOR COMMUNICATING ARTERY
C2882303|T047|I60.31|ICD10CM|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM RIGHT POSTERIOR COMMUNICATING ARTERY|NTRM SUBARACH HEMOR FROM RIGHT POST COMMUNICATING ARTERY
C2882302|T047|I60.30|ICD10CM|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM UNSPECIFIED POSTERIOR COMMUNICATING ARTERY|NTRM SUBARACH HEMOR FROM UNSP POSTERIOR COMMUNICATING ARTERY
C2833952|T037|S14.129D|ICD10CM|CENTRAL CORD SYNDROME AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|CENTRAL CORD SYND AT UNSP LEVEL OF CERV SPINAL CORD, SUBS
C2833951|T037|S14.129A|ICD10CM|CENTRAL CORD SYNDROME AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|CENTRAL CORD SYND AT UNSP LEVEL OF CERV SPINAL CORD, INIT
C2887447|T047|J44.1|ICD10CM|CHRONIC OBSTRUCTIVE PULMONARY DISEASE WITH (ACUTE) EXACERBATION|DECOMPENSATED COPD WITH (ACUTE) EXACERBATION
C2855940|T037|S68.128S|ICD10CM|PARTIAL TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF OTHER FINGER, SEQUELA|PARTIAL TRAUMATIC MCP AMPUTATION OF FINGER, SEQUELA
C4269382|T037|S02.40AS|ICD10CM|MALAR FRACTURE, RIGHT SIDE, SEQUELA|MALAR FRACTURE, RIGHT SIDE, SEQUELA
C4270348|T046|T83.598A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO OTHER PROSTHETIC DEVICE, IMPLANT AND GRAFT IN URINARY SYSTEM, INITIAL ENCOUNTER|I/I REACT D/T OTHER PROSTH DEV/GRFT URN SYS, INIT
C2876141|T037|T31.44|ICD10CM|BURNS INVOLVING 40-49% OF BODY SURFACE WITH 40-49% THIRD DEGREE BURNS|BURNS OF 40-49% OF BODY SURFACE W 40-49% THIRD DEGREE BURNS
C2876138|T037|T31.41|ICD10CM|BURNS INVOLVING 40-49% OF BODY SURFACE WITH 10-19% THIRD DEGREE BURNS|BURNS OF 40-49% OF BODY SURFACE W 10-19% THIRD DEGREE BURNS
C2876140|T037|T31.43|ICD10CM|BURNS INVOLVING 40-49% OF BODY SURFACE WITH 30-39% THIRD DEGREE BURNS|BURNS OF 40-49% OF BODY SURFACE W 30-39% THIRD DEGREE BURNS
C2876139|T037|T31.42|ICD10CM|BURNS INVOLVING 40-49% OF BODY SURFACE WITH 20-29% THIRD DEGREE BURNS|BURNS OF 40-49% OF BODY SURFACE W 20-29% THIRD DEGREE BURNS
C2890445|T037|T84.028A|ICD10CM|DISLOCATION OF OTHER INTERNAL JOINT PROSTHESIS, INITIAL ENCOUNTER|DISLOCATION OF OTHER INTERNAL JOINT PROSTHESIS, INIT ENCNTR
C2891342|T037|T87.9|ICD10CM|UNSPECIFIED COMPLICATIONS OF AMPUTATION STUMP|UNSPECIFIED COMPLICATIONS OF AMPUTATION STUMP
C2838214|T037|S32.456A|ICD10CM|NONDISPLACED TRANSVERSE FRACTURE OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED TRANSVERSE FRACTURE OF UNSP ACETABULUM, INIT
C2858028|T037|S72.351A|ICD10CM|DISPLACED COMMINUTED FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED COMMINUTED FRACTURE OF SHAFT OF RIGHT FEMUR, INIT
C2858029|T037|S72.351B|ICD10CM|DISPLACED COMMINUTED FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL COMMNT FX SHAFT OF R FEMUR, INIT FOR OPN FX TYPE I/2
C2858030|T037|S72.351C|ICD10CM|DISPLACED COMMINUTED FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL COMMNT FX SHAFT OF R FEMR, INIT FOR OPN FX TYPE 3A/B/C
C2887413|T047|J14|ICD10CM|PNEUMONIA DUE TO HEMOPHILUS INFLUENZAE|BRONCHOPNEUMONIA DUE TO H. INFLUENZAE
C2887412|T047|J13|ICD10CM|PNEUMONIA DUE TO STREPTOCOCCUS PNEUMONIAE|BRONCHOPNEUMONIA DUE TO S. PNEUMONIAE
C2887784|T047|K50.914|ICD10CM|CROHN'S DISEASE, UNSPECIFIED, WITH ABSCESS|CROHN'S DISEASE, UNSPECIFIED, WITH ABSCESS
C2888935|T047|M01.X29|ICD10CM|DIRECT INFECTION OF UNSPECIFIED ELBOW IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIR INFCT OF UNSP ELBOW IN INFEC/PARASTC DIS CLASSD ELSWHR
C2887782|T047|K50.912|ICD10CM|CROHN'S DISEASE, UNSPECIFIED, WITH INTESTINAL OBSTRUCTION|CROHN'S DISEASE, UNSPECIFIED, WITH INTESTINAL OBSTRUCTION
C2887783|T047|K50.913|ICD10CM|CROHN'S DISEASE, UNSPECIFIED, WITH FISTULA|CROHN'S DISEASE, UNSPECIFIED, WITH FISTULA
C2838215|T037|S32.456B|ICD10CM|NONDISPLACED TRANSVERSE FRACTURE OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP TRANSVERSE FX UNSP ACETABULUM, INIT FOR OPN FX
C2905748|T037|X77.9XXS|ICD10CM|INTENTIONAL SELF-HARM BY UNSPECIFIED HOT OBJECTS, SEQUELA|INTENTIONAL SELF-HARM BY UNSPECIFIED HOT OBJECTS, SEQUELA
C2887785|T047|K50.918|ICD10CM|CROHN'S DISEASE, UNSPECIFIED, WITH OTHER COMPLICATION|CROHN'S DISEASE, UNSPECIFIED, WITH OTHER COMPLICATION
C2888933|T047|M01.X21|ICD10CM|DIRECT INFECTION OF RIGHT ELBOW IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIRECT INFCT OF R ELBOW IN INFEC/PARASTC DIS CLASSD ELSWHR
C2888934|T047|M01.X22|ICD10CM|DIRECT INFECTION OF LEFT ELBOW IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIRECT INFCT OF L ELBOW IN INFEC/PARASTC DIS CLASSD ELSWHR
C2905746|T037|X77.9XXA|ICD10CM|INTENTIONAL SELF-HARM BY UNSPECIFIED HOT OBJECTS, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY UNSP HOT OBJECTS, INIT ENCNTR
C2905747|T037|X77.9XXD|ICD10CM|INTENTIONAL SELF-HARM BY UNSPECIFIED HOT OBJECTS, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY UNSP HOT OBJECTS, SUBS ENCNTR
C2901349|T046|M84.576A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, UNSPECIFIED FOOT, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, UNSP FOOT, INIT
C4270603|T046|T85.738A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO OTHER NERVOUS SYSTEM DEVICE, IMPLANT OR GRAFT, INITIAL ENCOUNTER|I/I REACT D/T OTHER NRV SYS DEVICE, IMPLNT OR GRAFT, INIT
C4268692|T047|M04.2|ICD10CM|CRYOPYRIN-ASSOCIATED PERIODIC SYNDROMES|NEONATAL ONSET MULTISYSTEMIC INFLAMMATORY DISORDER [NOMID]
C4268691|T047|M04.1|ICD10CM|PERIODIC FEVER SYNDROMES|TUMOR NECROSIS FACTOR RECEPTOR ASSOCIATED PERIODIC SYNDROME [TRAPS]
C2882964|T047|I70.669|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, UNSPECIFIED EXTREMITY|ATHSCL NONBIOL BYPASS OF THE EXTRM W GANGRENE, UNSP EXTRM
C4268696|T047|M04.9|ICD10CM|AUTOINFLAMMATORY SYNDROME, UNSPECIFIED|AUTOINFLAMMATORY SYNDROME, UNSPECIFIED
C4268694|T047|M04.8|ICD10CM|OTHER AUTOINFLAMMATORY SYNDROMES|PERIODIC FEVER, APHTHOUS STOMATITIS, PHARYNGITIS, AND ADENOPATHY SYNDROME [PFAPA]
C2902029|T046|M87.178|ICD10CM|OSTEONECROSIS DUE TO DRUGS, LEFT TOE(S)|OSTEONECROSIS DUE TO DRUGS, LEFT TOE(S)
C2902030|T046|M87.179|ICD10CM|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED TOE(S)|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED TOE(S)
C2902022|T046|M87.171|ICD10CM|OSTEONECROSIS DUE TO DRUGS, RIGHT ANKLE|OSTEONECROSIS DUE TO DRUGS, RIGHT ANKLE
C2902023|T046|M87.172|ICD10CM|OSTEONECROSIS DUE TO DRUGS, LEFT ANKLE|OSTEONECROSIS DUE TO DRUGS, LEFT ANKLE
C2902024|T046|M87.173|ICD10CM|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED ANKLE|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED ANKLE
C2902025|T046|M87.174|ICD10CM|OSTEONECROSIS DUE TO DRUGS, RIGHT FOOT|OSTEONECROSIS DUE TO DRUGS, RIGHT FOOT
C2902026|T046|M87.175|ICD10CM|OSTEONECROSIS DUE TO DRUGS, LEFT FOOT|OSTEONECROSIS DUE TO DRUGS, LEFT FOOT
C2902027|T046|M87.176|ICD10CM|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED FOOT|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED FOOT
C2902028|T046|M87.177|ICD10CM|OSTEONECROSIS DUE TO DRUGS, RIGHT TOE(S)|OSTEONECROSIS DUE TO DRUGS, RIGHT TOE(S)
C4267981|T047|E09.3519|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|DRUG/CHEM DIAB WITH PROLIF DIAB RTNOP WITH MCLR EDEMA, UNSP
C0019034|T047|D57.2|ICD10CM|SICKLE-CELL/HB-C DISEASE WITHOUT CRISIS|HB-S/HB-C DISEASE
C2070032|T046||ICD10CM|VITREOUS HEMORRHAGE, RIGHT EYE
C2887311|T047|I87.332|ICD10CM|CHRONIC VENOUS HYPERTENSION (IDIOPATHIC) WITH ULCER AND INFLAMMATION OF LEFT LOWER EXTREMITY|CHRONIC VENOUS HTN W ULCER AND INFLAMMATION OF L LOW EXTREM
C2881056|T046|H43.13|ICD10CM|VITREOUS HEMORRHAGE, BILATERAL|VITREOUS HEMORRHAGE, BILATERAL
C2070033|T046||ICD10CM|VITREOUS HEMORRHAGE, LEFT EYE
C4267978|T047|E09.3511|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|DRUG/CHEM DIAB WITH PROLIF DIAB RTNOP WITH MCLR EDEMA, R EYE
C4267979|T047|E09.3512|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|DRUG/CHEM DIAB WITH PROLIF DIAB RTNOP WITH MCLR EDEMA, L EYE
C4267916|T047|E08.3419|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|DIABETES WITH SEVERE NONP RTNOP WITH MACULAR EDEMA, UNSP
C2858661|T037|S72.442A|ICD10CM|DISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF LOWER EPIPHYSIS (SEPARATION) OF LEFT FEMUR, INIT
C2858663|T037|S72.442C|ICD10CM|DISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF LOW EPIPHY (SEPARATION) OF L FEMR, 7THC
C2858662|T037|S72.442B|ICD10CM|DISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF LOW EPIPHY (SEPARATION) OF L FEMR, 7THB
C2889102|T047|M02.872|ICD10CM|OTHER REACTIVE ARTHROPATHIES, LEFT ANKLE AND FOOT|OTHER REACTIVE ARTHROPATHIES, LEFT ANKLE AND FOOT
C2889101|T047|M02.871|ICD10CM|OTHER REACTIVE ARTHROPATHIES, RIGHT ANKLE AND FOOT|OTHER REACTIVE ARTHROPATHIES, RIGHT ANKLE AND FOOT
C2882960|T047|I70.661|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, RIGHT LEG|ATHSCL NONBIOL BYPASS OF THE EXTRM W GANGRENE, RIGHT LEG
C2837714|T037|S32.122B|ICD10CM|SEVERELY DISPLACED ZONE II FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|SEVERELY DISPLACED ZONE II FX SACRUM, INIT FOR OPN FX
C2889103|T047|M02.879|ICD10CM|OTHER REACTIVE ARTHROPATHIES, UNSPECIFIED ANKLE AND FOOT|OTHER REACTIVE ARTHROPATHIES, UNSPECIFIED ANKLE AND FOOT
C2838658|T037|S34.115D|ICD10CM|COMPLETE LESION OF L5 LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION OF L5 LEVEL OF LUMBAR SPINAL CORD, SUBS
C2838657|T037|S34.115A|ICD10CM|COMPLETE LESION OF L5 LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION OF L5 LEVEL OF LUMBAR SPINAL CORD, INIT
C0014868|T047|K20|ICD10CM|ESOPHAGITIS, UNSPECIFIED|ESOPHAGITIS
C0375352|T047|K20.8|ICD10CM|OTHER ESOPHAGITIS|OTHER ESOPHAGITIS
C0341106|T047|K20.0|ICD10CM|EOSINOPHILIC ESOPHAGITIS|EOSINOPHILIC ESOPHAGITIS
C2889126|T047|M05.061|ICD10CM|FELTY'S SYNDROME, RIGHT KNEE|FELTY'S SYNDROME, RIGHT KNEE
C2889127|T047|M05.062|ICD10CM|FELTY'S SYNDROME, LEFT KNEE|FELTY'S SYNDROME, LEFT KNEE
C2838659|T037|S34.115S|ICD10CM|COMPLETE LESION OF L5 LEVEL OF LUMBAR SPINAL CORD, SEQUELA|COMPLETE LESION OF L5 LEVEL OF LUMBAR SPINAL CORD, SEQUELA
C2900511|T046|M80.852A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, LEFT FEMUR, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, LEFT FEMUR, INIT
C2842079|T191|C50.019|ICD10CM|MALIGNANT NEOPLASM OF NIPPLE AND AREOLA, UNSPECIFIED FEMALE BREAST|MALIGNANT NEOPLASM OF NIPPLE AND AREOLA, UNSP FEMALE BREAST
C3469323|T047|M05.069|ICD10CM|FELTY'S SYNDROME, UNSPECIFIED KNEE|FELTY'S SYNDROME, UNSPECIFIED KNEE
C2902865|T047|N01.9|ICD10CM|RAPIDLY PROGRESSIVE NEPHRITIC SYNDROME WITH UNSPECIFIED MORPHOLOGIC CHANGES|RAPIDLY PROGR NEPHRITIC SYNDROME W UNSP MORPHOLOGIC CHANGES
C2902864|T047|N01.8|ICD10CM|RAPIDLY PROGRESSIVE NEPHRITIC SYNDROME WITH OTHER MORPHOLOGIC CHANGES|RAPIDLY PROGR NEPHRITIC SYNDROME W OTH MORPHOLOGIC CHANGES
C2884980|T037|T59.892S|ICD10CM|TOXIC EFFECT OF OTHER SPECIFIED GASES, FUMES AND VAPORS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF GASES, FUMES AND VAPORS, SELF-HARM, SEQUELA
C2902859|T047|N01.1|ICD10CM|RAPIDLY PROGRESSIVE NEPHRITIC SYNDROME WITH FOCAL AND SEGMENTAL GLOMERULAR LESIONS|RAPIDLY PROGRESSIVE NEPHRITIC SYNDROME WITH FOCAL GLOMERULONEPHRITIS
C2902856|T047|N01.0|ICD10CM|RAPIDLY PROGRESSIVE NEPHRITIC SYNDROME WITH MINOR GLOMERULAR ABNORMALITY|RAPIDLY PROGRESSIVE NEPHRITIC SYNDROME WITH MINIMAL CHANGE LESION
C0451732|T047|N01.3|DMDICD10|RAPIDLY PROGRESSIVE NEPHRITIC SYNDROME WITH DIFFUSE MESANGIAL PROLIFERATIVE GLOMERULONEPHRITIS|RAPID-PROGRESSIVES NEPHRITISCHES SYNDROM: DIFFUSE MESANGIOPROLIFERATIVE GLOMERULONEPHRITIS
C0451731|T047|N01.2|DMDICD10|RAPIDLY PROGRESSIVE NEPHRITIC SYNDROME WITH DIFFUSE MEMBRANOUS GLOMERULONEPHRITIS|RAPID-PROGRESSIVES NEPHRITISCHES SYNDROM: DIFFUSE MEMBRANOESE GLOMERULONEPHRITIS
C2902860|T047|N01.5|ICD10CM|RAPIDLY PROGRESSIVE NEPHRITIC SYNDROME WITH DIFFUSE MESANGIOCAPILLARY GLOMERULONEPHRITIS|RAPIDLY PROGRESSIVE NEPHRITIC SYNDROME WITH MEMBRANOPROLIFERATIVE GLOMERULONEPHRITIS, TYPES 1 AND 3, OR NOS
C0451733|T047|N01.4|DMDICD10|RAPIDLY PROGRESSIVE NEPHRITIC SYNDROME WITH DIFFUSE ENDOCAPILLARY PROLIFERATIVE GLOMERULONEPHRITIS|RAPID-PROGRESSIVES NEPHRITISCHES SYNDROM: DIFFUSE ENDOKAPILLAER-PROLIFERATIVE GLOMERULONEPHRITIS
C2902862|T047|N01.7|ICD10CM|RAPIDLY PROGRESSIVE NEPHRITIC SYNDROME WITH DIFFUSE CRESCENTIC GLOMERULONEPHRITIS|RAPIDLY PROGRESSIVE NEPHRITIC SYNDROME WITH EXTRACAPILLARY GLOMERULONEPHRITIS
C2902861|T047|N01.6|ICD10CM|RAPIDLY PROGRESSIVE NEPHRITIC SYNDROME WITH DENSE DEPOSIT DISEASE|RAPIDLY PROGRESSIVE NEPHRITIC SYNDROME WITH MEMBRANOPROLIFERATIVE GLOMERULONEPHRITIS, TYPE 2
C0838482|T047||ICD10CM|ANKYLOSING SPONDYLITIS OF MULTIPLE SITES IN SPINE
C0838483|T047||ICD10CM|ANKYLOSING SPONDYLITIS OF OCCIPITO-ATLANTO-AXIAL REGION
C0838484|T047||ICD10CM|ANKYLOSING SPONDYLITIS OF CERVICAL REGION
C0838485|T047||ICD10CM|ANKYLOSING SPONDYLITIS OF CERVICOTHORACIC REGION
C0838486|T047||ICD10CM|ANKYLOSING SPONDYLITIS OF THORACIC REGION
C0838487|T047||ICD10CM|ANKYLOSING SPONDYLITIS OF THORACOLUMBAR REGION
C0838488|T047||ICD10CM|ANKYLOSING SPONDYLITIS LUMBAR REGION
C0838489|T047||ICD10CM|ANKYLOSING SPONDYLITIS OF LUMBOSACRAL REGION
C0838490|T047||ICD10CM|ANKYLOSING SPONDYLITIS SACRAL AND SACROCOCCYGEAL REGION
C2895253|T047|M45.9|ICD10CM|ANKYLOSING SPONDYLITIS OF UNSPECIFIED SITES IN SPINE|ANKYLOSING SPONDYLITIS OF UNSPECIFIED SITES IN SPINE
C2879747|T037|T47.3X2A|ICD10CM|POISONING BY SALINE AND OSMOTIC LAXATIVES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY SALINE AND OSMOTIC LAXATIVES, SELF-HARM, INIT
C2977715|T037|S02.609S|ICD10CM|FRACTURE OF MANDIBLE, UNSPECIFIED, SEQUELA|FRACTURE OF MANDIBLE, UNSPECIFIED, SEQUELA
C2838495|T037|S32.810A|ICD10CM|MULTIPLE FRACTURES OF PELVIS WITH STABLE DISRUPTION OF PELVIC RING, INITIAL ENCOUNTER FOR CLOSED FRACTURE|MULTIPLE FX OF PELVIS W STABLE DISRUPT OF PELVIC RING, INIT
C2893631|T047|M12.019|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], UNSPECIFIED SHOULDER|CHRONIC POSTRHEUMATIC ARTHROPATHY, UNSPECIFIED SHOULDER
C4267911|T047|E08.3393|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|DIABETES WITH MODERATE NONP RTNOP WITHOUT MACULAR EDEMA, BI
C4267910|T047|E08.3392|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|DIAB WITH MODERATE NONP RTNOP WITHOUT MACULAR EDEMA, L EYE
C4267909|T047|E08.3391|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|DIAB WITH MODERATE NONP RTNOP WITHOUT MACULAR EDEMA, R EYE
C4267912|T047|E08.3399|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|DIAB WITH MODERATE NONP RTNOP WITHOUT MACULAR EDEMA, UNSP
C2890467|T037|T84.033A|ICD10CM|MECHANICAL LOOSENING OF INTERNAL LEFT KNEE PROSTHETIC JOINT, INITIAL ENCOUNTER|MECH LOOSENING OF INTERNAL LEFT KNEE PROSTHETIC JOINT, INIT
C2848421|T037|S58.112S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN ELBOW AND WRIST, LEFT ARM, SEQUELA|COMPLETE TRAUM AMP AT LEV BETW ELBOW AND WRS, LEFT ARM, SQLA
C2879000|T037|T44.992A|ICD10CM|POISONING BY OTHER DRUG PRIMARILY AFFECTING THE AUTONOMIC NERVOUS SYSTEM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY OTH DRUG AFF THE AUTONM NERVOUS SYS, SLF-HRM, INIT
C2902130|T046|M87.822|ICD10CM|OTHER OSTEONECROSIS, LEFT HUMERUS|OTHER OSTEONECROSIS, LEFT HUMERUS
C2902129|T046|M87.821|ICD10CM|OTHER OSTEONECROSIS, RIGHT HUMERUS|OTHER OSTEONECROSIS, RIGHT HUMERUS
C2879002|T037|T44.992S|ICD10CM|POISONING BY OTHER DRUG PRIMARILY AFFECTING THE AUTONOMIC NERVOUS SYSTEM, INTENTIONAL SELF-HARM, SEQUELA|POISN BY OTH DRUG AFF THE AUTONM NRV SYS, SLF-HRM, SEQUELA
C2833591|T037|S12.601A|ICD10CM|UNSPECIFIED NONDISPLACED FRACTURE OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP NONDISP FX OF SEVENTH CERVICAL VERTEBRA, INIT
C2833592|T037|S12.601B|ICD10CM|UNSPECIFIED NONDISPLACED FRACTURE OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP NONDISP FX OF SEVENTH CERVCAL VERTEBRA, INIT FOR OPN FX
C2902131|T046|M87.82|ICD10CM|OTHER OSTEONECROSIS, UNSPECIFIED HUMERUS|OTHER OSTEONECROSIS, HUMERUS
C2835858|T037|S24.159D|ICD10CM|OTHER INCOMPLETE LESION AT UNSPECIFIED LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|OTH INCMPL LESION AT UNSP LEVEL OF THOR SPINAL CORD, SUBS
C4237013|T048|F15.980|ICD10CM|OTHER STIMULANT USE, UNSPECIFIED WITH STIMULANT-INDUCED ANXIETY DISORDER|CAFFEINE INDUCED ANXIETY DISORDER, WITHOUT USE DISORDER
C2838712|T037|S34.3XXA|ICD10CM|INJURY OF CAUDA EQUINA, INITIAL ENCOUNTER|INJURY OF CAUDA EQUINA, INITIAL ENCOUNTER
C2832036|T037|S06.2X6A|ICD10CM|DIFFUSE TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|DIFFUSE TBI W LOC >24 HR W/O RET CONSC W SURV, INIT
C2902437|T047|M90.541|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, RIGHT HAND|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, RIGHT HAND
C2875112|T047|G40.401|ICD10CM|OTHER GENERALIZED EPILEPSY AND EPILEPTIC SYNDROMES, NOT INTRACTABLE, WITH STATUS EPILEPTICUS|OTH GENERALIZED EPILEPSY, NOT INTRACTABLE, W STAT EPI
C0524851|T047|G31.9|DMDICD10|DEGENERATIVE DISEASE OF NERVOUS SYSTEM, UNSPECIFIED|DEGENERATIVE KRANKHEIT DES NERVENSYSTEMS, NICHT NAEHER BEZEICHNET
C2875113|T047|G40.409|ICD10CM|OTHER GENERALIZED EPILEPSY AND EPILEPTIC SYNDROMES, NOT INTRACTABLE, WITHOUT STATUS EPILEPTICUS|OTH GENERALIZED EPILEPSY, NOT INTRACTABLE, W/O STAT EPI
C0494465|T047|G31.1|DMDICD10|SENILE DEGENERATION OF BRAIN, NOT ELSEWHERE CLASSIFIED|SENILE DEGENERATION DES GEHIRNS, ANDERENORTS NICHT KLASSIFIZIERT
C2832038|T037|S06.2X6S|ICD10CM|DIFFUSE TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|DIFFUSE TBI W LOC >24 HR W/O RET CONSC W SURV, SEQUELA
C2931917|T047|G31.2|ICD10CM|DEGENERATION OF NERVOUS SYSTEM DUE TO ALCOHOL|ALCOHOLIC ENCEPHALOPATHY
C2900569|T046|M80.88XA|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, VERTEBRA(E), INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, VERTEBRA(E), INIT
C2890122|T037|T82.598A|ICD10CM|OTHER MECHANICAL COMPLICATION OF OTHER CARDIAC AND VASCULAR DEVICES AND IMPLANTS, INITIAL ENCOUNTER|MECH COMPL OF CARDIAC AND VASCULAR DEVICES AND IMPLNT, INIT
C2882191|T047|I25.738|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL CORONARY ARTERY BYPASS GRAFT(S) WITH OTHER FORMS OF ANGINA PECTORIS|ATHSCL NONAUTOLOGOUS BIOLOGICAL CABG W OTH ANGINA PECTORIS
C2882192|T047|I25.739|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL CORONARY ARTERY BYPASS GRAFT(S) WITH UNSPECIFIED ANGINA PECTORIS|ATHSCL NONAUTOLOGOUS BIOLOGICAL CABG W UNSP ANGINA PECTORIS
C2882189|T047|I25.730|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL CORONARY ARTERY BYPASS GRAFT(S) WITH UNSTABLE ANGINA PECTORIS|ATHSCL NONAUTOLOGOUS BIOLOGICAL CABG W UNSTABLE ANG PCTRS
C2882190|T047|I25.731|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL CORONARY ARTERY BYPASS GRAFT(S) WITH ANGINA PECTORIS WITH DOCUMENTED SPASM|ATHSCL NONAUT BIOLOGICAL CABG W ANG PCTRS W DOCUMENTED SPASM
C2838143|T037|S32.442A|ICD10CM|DISPLACED FRACTURE OF POSTERIOR COLUMN [ILIOISCHIAL] OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF POSTERIOR COLUMN OF LEFT ACETABULUM, INIT
C2838144|T037|S32.442B|ICD10CM|DISPLACED FRACTURE OF POSTERIOR COLUMN [ILIOISCHIAL] OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISP FX OF POSTERIOR COLUMN OF LEFT ACETAB, INIT FOR OPN FX
C2833866|T037|S14.106A|ICD10CM|UNSPECIFIED INJURY AT C6 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY AT C6 LEVEL OF CERVICAL SPINAL CORD, INIT ENCNTR
C4267933|T047|E08.3533|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, BILATERAL|DIAB WITH PROLIF DIABETIC RTNOP WITH TRCTN DTCH N-MCLA, BI
C4267932|T047|E08.3532|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, LEFT EYE|DIAB WITH PROLIF DIAB RTNOP WITH TRCTN DTCH N-MCLA, LEFT EYE
C4267931|T047|E08.3531|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, RIGHT EYE|DIAB WITH PROLIF DIAB RTNOP WITH TRCTN DTCH N-MCLA, R EYE
C2885458|T037|T63.112A|ICD10CM|TOXIC EFFECT OF VENOM OF GILA MONSTER, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF GILA MONSTER, SELF-HARM, INIT
C2837532|T037|S32.022B|ICD10CM|UNSTABLE BURST FRACTURE OF SECOND LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSTABLE BURST FX SECOND LUM VERTEBRA, INIT FOR OPN FX
C4267934|T047|E08.3539|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, UNSPECIFIED EYE|DIAB WITH PROLIF DIABETIC RTNOP WITH TRCTN DTCH N-MCLA, UNSP
C2853983|T191|C84.73|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-NEGATIVE, INTRA-ABDOMINAL LYMPH NODES|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-NEG, INTRA-ABD NODES
C2853982|T191|C84.72|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-NEGATIVE, INTRATHORACIC LYMPH NODES|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-NEG, INTRATHORAC NODES
C2853981|T191|C84.71|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-NEGATIVE, LYMPH NODES OF HEAD, FACE, AND NECK|ANAPLSTC LG CELL LYMPH, ALK-NEG, NODES OF HEAD, FACE, AND NK
C2853980|T191|C84.70|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-NEGATIVE, UNSPECIFIED SITE|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-NEGATIVE, UNSP SITE
C2853987|T191||ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-NEGATIVE, SPLEEN
C2853986|T191|C84.76|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-NEGATIVE, INTRAPELVIC LYMPH NODES|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-NEG, INTRAPELV NODES
C2853985|T191|C84.75|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-NEGATIVE, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|ANAPLSTC LG CELL LYMPH, ALK-NEG, NODES OF ING RGN & LOW LMB
C2853984|T191|C84.74|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-NEGATIVE, LYMPH NODES OF AXILLA AND UPPER LIMB|ANAPLSTC LG CELL LYMPH, ALK-NEG, NODES OF AXLA AND UPR LIMB
C2853989|T191|C84.79|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-NEGATIVE, EXTRANODAL AND SOLID ORGAN SITES|ANAPLSTC LG CELL LYMPH, ALK-NEG, EXTRNOD AND SOLID ORG SITES
C2853988|T191|C84.78|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-NEGATIVE, LYMPH NODES OF MULTIPLE SITES|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-NEG, NODES MULT SITE
C2833279|T037|S12.14XB|ICD10CM|TYPE III TRAUMATIC SPONDYLOLISTHESIS OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE III TRAUM SPONDYLOLYSIS OF 2ND CERVCAL VERT, 7THB
C2833278|T037|S12.14XA|ICD10CM|TYPE III TRAUMATIC SPONDYLOLISTHESIS OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE III TRAUM SPONDYLOLYSIS OF SECOND CERVCAL VERT, INIT
C2888796|T047|M00.012|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, LEFT SHOULDER|STAPHYLOCOCCAL ARTHRITIS, LEFT SHOULDER
C2910373|T049|Q93.89|ICD10CM|OTHER DELETIONS FROM THE AUTOSOMES|DELETIONS IDENTIFIED BY IN SITU HYBRIDIZATION (ISH)
C2888795|T047|M00.011|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, RIGHT SHOULDER|STAPHYLOCOCCAL ARTHRITIS, RIGHT SHOULDER
C2856691|T037|S72.031B|ICD10CM|DISPLACED MIDCERVICAL FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPLACED MIDCERVICAL FX R FEMUR, INIT FOR OPN FX TYPE I/2
C2886035|T037|T65.222S|ICD10CM|TOXIC EFFECT OF TOBACCO CIGARETTES, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF TOBACCO CIGARETTES, SELF-HARM, SEQUELA
C0220704|T047|Q93.81|ICD10CM|VELO-CARDIO-FACIAL SYNDROME|DELETION 22Q11.2
C2888797|T047|M00.019|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, UNSPECIFIED SHOULDER|STAPHYLOCOCCAL ARTHRITIS, UNSPECIFIED SHOULDER
C2861598|T191||ICD10CM|ACUTE MYELOMONOCYTIC LEUKEMIA, NOT HAVING ACHIEVED REMISSION
C0836973|T191||ICD10AM|ACUTE MYELOMONOCYTIC LEUKEMIA, IN REMISSION
C2861599|T191||ICD10CM|ACUTE MYELOMONOCYTIC LEUKEMIA, IN RELAPSE
C2882812|T047|I70.419|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, UNSPECIFIED EXTREMITY|ATHSCL AUTOL VEIN BYPASS OF EXTRM W INTRMT CLAUD, UNSP EXTRM
C2882811|T047|I70.418|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, OTHER EXTREMITY|ATHSCL AUTOL VEIN BYPASS OF EXTRM W INTRMT CLAUD, OTH EXTRM
C2882222|T047|I26.99|ICD10CM|OTHER PULMONARY EMBOLISM WITHOUT ACUTE COR PULMONALE|OTHER PULMONARY EMBOLISM WITHOUT ACUTE COR PULMONALE
C2882808|T047|I70.411|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, RIGHT LEG|ATHSCL AUTOL VEIN BYPASS OF EXTRM W INTRMT CLAUD, RIGHT LEG
C3264367|T047|I26.92|ICD10CM|SADDLE EMBOLUS OF PULMONARY ARTERY WITHOUT ACUTE COR PULMONALE|SADDLE EMBOLUS OF PULMONARY ARTERY W/O ACUTE COR PULMONALE
C2882810|T047|I70.413|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, BILATERAL LEGS|ATHSCL AUTOL VEIN BYPASS OF EXTRM W INTRMT CLAUD, BI LEGS
C2882220|T047|I26.90|ICD10CM|SEPTIC PULMONARY EMBOLISM WITHOUT ACUTE COR PULMONALE|SEPTIC PULMONARY EMBOLISM WITHOUT ACUTE COR PULMONALE
C2835298|T037|S22.040A|ICD10CM|WEDGE COMPRESSION FRACTURE OF FOURTH THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|WEDGE COMPRESSION FRACTURE OF FOURTH THORACIC VERTEBRA, INIT
C2835299|T037|S22.040B|ICD10CM|WEDGE COMPRESSION FRACTURE OF FOURTH THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|WEDGE COMPRSN FX FOURTH THOR VERTEBRA, INIT FOR OPN FX
C2905721|T037|X75.XXXS|ICD10CM|INTENTIONAL SELF-HARM BY EXPLOSIVE MATERIAL, SEQUELA|INTENTIONAL SELF-HARM BY EXPLOSIVE MATERIAL, SEQUELA
C0178416|T047||ICD10CM|APLASTIC ANEMIA, UNSPECIFIED
C4267948|T047|E08.3599|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|DIAB WITH PROLIF DIABETIC RTNOP WITHOUT MACULAR EDEMA, UNSP
C2842123|T191|C50.621|ICD10CM|MALIGNANT NEOPLASM OF AXILLARY TAIL OF RIGHT MALE BREAST|MALIGNANT NEOPLASM OF AXILLARY TAIL OF RIGHT MALE BREAST
C0271909|T047|D61.1|DMDICD10|DRUG-INDUCED APLASTIC ANEMIA|ARZNEIMITTELINDUZIERTE APLASTISCHE ANAEMIE
C0348890|T047|D61.3|DMDICD10|IDIOPATHIC APLASTIC ANEMIA|IDIOPATHISCHE APLASTISCHE ANAEMIE
C0494236|T047|D61.2|DMDICD10|APLASTIC ANEMIA DUE TO OTHER EXTERNAL AGENTS|APLASTISCHE ANAEMIE INFOLGE SONSTIGER AEUSSERER URSACHEN
C2902381|T047|M89.679|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, UNSPECIFIED ANKLE AND FOOT|OSTEOPATHY AFTER POLIOMYELITIS, UNSPECIFIED ANKLE AND FOOT
C2853995|T191|C84.94|ICD10CM|MATURE T/NK-CELL LYMPHOMAS, UNSPECIFIED, LYMPH NODES OF AXILLA AND UPPER LIMB|MATURE T/NK-CELL LYMPH, UNSP, NODES OF AXILLA AND UPPER LIMB
C2901813|T047|M86.161|ICD10CM|OTHER ACUTE OSTEOMYELITIS, RIGHT TIBIA AND FIBULA|OTHER ACUTE OSTEOMYELITIS, RIGHT TIBIA AND FIBULA
C2901814|T047|M86.162|ICD10CM|OTHER ACUTE OSTEOMYELITIS, LEFT TIBIA AND FIBULA|OTHER ACUTE OSTEOMYELITIS, LEFT TIBIA AND FIBULA
C2879466|T037|T46.3X2A|ICD10CM|POISONING BY CORONARY VASODILATORS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY CORONARY VASODILATORS, SELF-HARM, INIT
C2887149|T047|I82.B12|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF LEFT SUBCLAVIAN VEIN|ACUTE EMBOLISM AND THROMBOSIS OF LEFT SUBCLAVIAN VEIN
C2843282|T037|S48.021A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT RIGHT SHOULDER JOINT, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION AT RIGHT SHOULDER JOINT, INIT
C2901815|T047|M86.169|ICD10CM|OTHER ACUTE OSTEOMYELITIS, UNSPECIFIED TIBIA AND FIBULA|OTHER ACUTE OSTEOMYELITIS, UNSPECIFIED TIBIA AND FIBULA
C2833287|T037|S12.150B|ICD10CM|OTHER TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH TRAUM DISPL SPONDYLOLYSIS OF 2ND CERVCAL VERT, 7THB
C4268476|T047|I63.033|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF BILATERAL CAROTID ARTERIES|CEREBRAL INFRC DUE TO THOMBOS OF BILATERAL CAROTID ARTERIES
C2882337|T047|I63.032|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF LEFT CAROTID ARTERY|CEREBRAL INFARCTION DUE TO THROMBOSIS OF LEFT CAROTID ARTERY
C2882336|T047|I63.031|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF RIGHT CAROTID ARTERY|CEREBRAL INFRC DUE TO THROMBOSIS OF RIGHT CAROTID ARTERY
C2879468|T037|T46.3X2S|ICD10CM|POISONING BY CORONARY VASODILATORS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY CORONARY VASODILATORS, SELF-HARM, SEQUELA
C2882338|T047|I63.039|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF UNSPECIFIED CAROTID ARTERY|CEREBRAL INFARCTION DUE TO THROMBOSIS OF UNSP CAROTID ARTERY
C2843284|T037|S48.021S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT RIGHT SHOULDER JOINT, SEQUELA|PARTIAL TRAUMATIC AMPUTATION AT R SHOULDER JT, SEQUELA
C2885626|T037|T63.422A|ICD10CM|TOXIC EFFECT OF VENOM OF ANTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF ANTS, INTENTIONAL SELF-HARM, INIT
C2889269|T047|M05.521|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT ELBOW|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT ELBOW
C2857413|T037|S72.134C|ICD10CM|NONDISPLACED APOPHYSEAL FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP APOPHYSEAL FX R FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2859144|T037|S73.002A|ICD10CM|UNSPECIFIED SUBLUXATION OF LEFT HIP, INITIAL ENCOUNTER|UNSPECIFIED SUBLUXATION OF LEFT HIP, INITIAL ENCOUNTER
C2889270|T047|M05.522|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT ELBOW|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2859181|T037|S73.016A|ICD10CM|POSTERIOR DISLOCATION OF UNSPECIFIED HIP, INITIAL ENCOUNTER|POSTERIOR DISLOCATION OF UNSPECIFIED HIP, INITIAL ENCOUNTER
C2834014|T037|S14.146D|ICD10CM|BROWN-SEQUARD SYNDROME AT C6 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|BROWN-SEQUARD SYNDROME AT C6, SUBS
C2889271|T047|M05.52|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF ELBOW
C2858423|T037|S72.416A|ICD10CM|NONDISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP UNSP CONDYLE FX LOWER END OF UNSP FEMUR, INIT
C2858424|T037|S72.416B|ICD10CM|NONDISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP UNSP CONDYLE FX LOW END UNSP FEMR, 7THB
C2858425|T037|S72.416C|ICD10CM|NONDISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP UNSP CONDYLE FX LOW END UNSP FEMR, 7THC
C2834015|T037|S14.146S|ICD10CM|BROWN-SEQUARD SYNDROME AT C6 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|BROWN-SEQUARD SYNDROME AT C6, SEQUELA
C2879975|T037|T48.202S|ICD10CM|POISONING BY UNSPECIFIED DRUGS ACTING ON MUSCLES, INTENTIONAL SELF-HARM, SEQUELA|POISN BY UNSP DRUGS ACTING ON MUSCLES, SELF-HARM, SEQUELA
C2889633|T047|M08.929|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, UNSPECIFIED ELBOW|JUVENILE ARTHRITIS, UNSPECIFIED, UNSPECIFIED ELBOW
C2889632|T047|M08.922|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, LEFT ELBOW|JUVENILE ARTHRITIS, UNSPECIFIED, LEFT ELBOW
C2889631|T047|M08.921|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, RIGHT ELBOW|JUVENILE ARTHRITIS, UNSPECIFIED, RIGHT ELBOW
C2889384|T047|M05.89|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF MULTIPLE SITES|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR MULT SITE
C2835850|T037|S24.153D|ICD10CM|OTHER INCOMPLETE LESION AT T7-T10 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|OTH INCOMPLETE LESION AT T7-T10, SUBS
C2835849|T037|S24.153A|ICD10CM|OTHER INCOMPLETE LESION AT T7-T10 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|OTH INCOMPLETE LESION AT T7-T10, INIT
C2889356|T047|M05.8|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED SITE|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR
C2879181|T037|T45.522S|ICD10CM|POISONING BY ANTITHROMBOTIC DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ANTITHROMBOTIC DRUGS, SELF-HARM, SEQUELA
C2873983|T047|E09.40|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH NEUROLOGICAL COMPLICATIONS WITH DIABETIC NEUROPATHY, UNSPECIFIED|DRUG/CHEM DIABETES W NEURO COMP W DIABETIC NEUROPATHY, UNSP
C2856588|T037|S72.021C|ICD10CM|DISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF EPIPHY (SEPARATION) (UPPER) OF R FEMR, 7THC
C2890846|T037|T84.614A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL FIXATION DEVICE OF RIGHT ULNA, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INT FIX OF RIGHT ULNA, INIT
C2879179|T037|T45.522A|ICD10CM|POISONING BY ANTITHROMBOTIC DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ANTITHROMBOTIC DRUGS, SELF-HARM, INIT
C2835851|T037|S24.153S|ICD10CM|OTHER INCOMPLETE LESION AT T7-T10 LEVEL OF THORACIC SPINAL CORD, SEQUELA|OTH INCOMPLETE LESION AT T7-T10, SEQUELA
C2879946|T037|T48.1X2A|ICD10CM|POISONING BY SKELETAL MUSCLE RELAXANTS [NEUROMUSCULAR BLOCKING AGENTS], INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY SKELETAL MUSCLE RELAXANTS, SELF-HARM, INIT
C4269361|T037|S02.400S|ICD10CM|MALAR FRACTURE, UNSPECIFIED SIDE, SEQUELA|MALAR FRACTURE, UNSPECIFIED SIDE, SEQUELA
C2895315|T037|M48.51XA|ICD10CM|COLLAPSED VERTEBRA, NOT ELSEWHERE CLASSIFIED, OCCIPITO-ATLANTO-AXIAL REGION, INITIAL ENCOUNTER FOR FRACTURE|COLLAPSED VERTEBRA, NEC, OCCIPITO-ATLANTO-AXIAL REGION, INIT
C2878146|T037|T42.4X2A|ICD10CM|POISONING BY BENZODIAZEPINES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY BENZODIAZEPINES, INTENTIONAL SELF-HARM, INIT
C0039145|T047|G95.0|DMDICD10|SYRINGOMYELIA AND SYRINGOBULBIA|SYRINGOMYELIE UND SYRINGOBULBIE
C0037928|T047|G95.9|DMDICD10|DISEASE OF SPINAL CORD, UNSPECIFIED|KRANKHEIT DES RUECKENMARKES, NICHT NAEHER BEZEICHNET
C4269357|T037|S02.400B|ICD10CM|MALAR FRACTURE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|MALAR FRACTURE, UNSPECIFIED SIDE, 7THB
C4269356|T037|S02.400A|ICD10CM|MALAR FRACTURE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|MALAR FRACTURE, UNSPECIFIED SIDE, INIT
C2878148|T037|T42.4X2S|ICD10CM|POISONING BY BENZODIAZEPINES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY BENZODIAZEPINES, INTENTIONAL SELF-HARM, SEQUELA
C2838029|T037|S32.414B|ICD10CM|NONDISPLACED FRACTURE OF ANTERIOR WALL OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP FX OF ANTERIOR WALL OF RIGHT ACETAB, INIT FOR OPN FX
C0149886|T047||ICD10CM|SIMPLE FEBRILE CONVULSIONS
C1719637|T047|R56.01|ICD10CM|COMPLEX FEBRILE CONVULSIONS|COMPLICATED FEBRILE SEIZURE
C2901581|T046|M84.676A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, UNSPECIFIED FOOT, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, UNSP FOOT, INIT FOR FX
C4267956|T047|E09.3213|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|DRUG/CHEM DIAB WITH MILD NONP RTNOP WITH MACULAR EDEMA, BI
C4267955|T047|E09.3212|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|DRUG/CHEM DIAB WITH MILD NONP RTNOP WITH MCLR EDEMA, L EYE
C4267954|T047|E09.3211|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|DRUG/CHEM DIAB WITH MILD NONP RTNOP WITH MCLR EDEMA, R EYE
C2856086|T037|S68.711A|ICD10CM|COMPLETE TRAUMATIC TRANSMETACARPAL AMPUTATION OF RIGHT HAND, INITIAL ENCOUNTER|COMPLETE TRAUMATIC TRANSMETCRPL AMP OF RIGHT HAND, INIT
C2838237|T037|S32.463B|ICD10CM|DISPLACED ASSOCIATED TRANSVERSE-POSTERIOR FRACTURE OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISPLACED ASSOC TRANSV/POST FX UNSP ACETAB, INIT FOR OPN FX
C0155733|T047|I70.0|DMDICD10|ATHEROSCLEROSIS OF AORTA|ATHEROSKLEROSE DER AORTA
C2882691|T047|I70.1|ICD10CM|ATHEROSCLEROSIS OF RENAL ARTERY|GOLDBLATT'S KIDNEY
C4267957|T047|E09.3219|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|DRUG/CHEM DIAB WITH MILD NONP RTNOP WITH MACULAR EDEMA, UNSP
C4268036|T047|E10.3512|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|TYPE 1 DIAB WITH PROLIF DIAB RTNOP WITH MACULAR EDEMA, L EYE
C4268037|T047|E10.3513|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|TYPE 1 DIAB WITH PROLIF DIAB RTNOP WITH MACULAR EDEMA, BI
C2835815|T037|S24.139S|ICD10CM|ANTERIOR CORD SYNDROME AT UNSPECIFIED LEVEL OF THORACIC SPINAL CORD, SEQUELA|ANT CORD SYNDROME AT UNSP LEVEL OF THOR SPINAL CORD, SEQUELA
C4268035|T047|E10.3511|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|TYPE 1 DIAB WITH PROLIF DIAB RTNOP WITH MACULAR EDEMA, R EYE
C2902103|T046|M87.346|ICD10CM|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED FINGER(S)|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED FINGER(S)
C2902102|T046|M87.345|ICD10CM|OTHER SECONDARY OSTEONECROSIS, LEFT FINGER(S)|OTHER SECONDARY OSTEONECROSIS, LEFT FINGER(S)
C4268038|T047|E10.3519|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|TYPE 1 DIAB WITH PROLIF DIAB RTNOP WITH MACULAR EDEMA, UNSP
C2902100|T046|M87.343|ICD10CM|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED HAND|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED HAND
C2902099|T046|M87.342|ICD10CM|OTHER SECONDARY OSTEONECROSIS, LEFT HAND|OTHER SECONDARY OSTEONECROSIS, LEFT HAND
C2902098|T046|M87.341|ICD10CM|OTHER SECONDARY OSTEONECROSIS, RIGHT HAND|OTHER SECONDARY OSTEONECROSIS, RIGHT HAND
C2835813|T037|S24.139A|ICD10CM|ANTERIOR CORD SYNDROME AT UNSPECIFIED LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|ANT CORD SYNDROME AT UNSP LEVEL OF THOR SPINAL CORD, INIT
C0023370|T047|I74.01|ICD10CM|SADDLE EMBOLUS OF ABDOMINAL AORTA|SADDLE EMBOLUS OF ABDOMINAL AORTA
C2835814|T037|S24.139D|ICD10CM|ANTERIOR CORD SYNDROME AT UNSPECIFIED LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|ANT CORD SYNDROME AT UNSP LEVEL OF THOR SPINAL CORD, SUBS
C3161092|T047|I74.09|ICD10CM|OTHER ARTERIAL EMBOLISM AND THROMBOSIS OF ABDOMINAL AORTA|OTHER ARTERIAL EMBOLISM AND THROMBOSIS OF ABDOMINAL AORTA
C2837853|T037|S32.315A|ICD10CM|NONDISPLACED AVULSION FRACTURE OF LEFT ILIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED AVULSION FRACTURE OF LEFT ILIUM, INIT
C2837854|T037|S32.315B|ICD10CM|NONDISPLACED AVULSION FRACTURE OF LEFT ILIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP AVULSION FRACTURE OF LEFT ILIUM, INIT FOR OPN FX
C2896530|T046|M80.031A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, RIGHT FOREARM, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, R FOREARM, INIT
C2885643|T037|T63.432A|ICD10CM|TOXIC EFFECT OF VENOM OF CATERPILLARS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF CATERPILLARS, SELF-HARM, INIT
C2885645|T037|T63.432S|ICD10CM|TOXIC EFFECT OF VENOM OF CATERPILLARS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF CATERPILLARS, SELF-HARM, SEQUELA
C2833487|T037|S12.450A|ICD10CM|OTHER TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH TRAUM DISPL SPONDYLOLYSIS OF FIFTH CERVCAL VERT, INIT
C2832060|T037|S06.301S|ICD10CM|UNSPECIFIED FOCAL TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|UNSP FOCAL TBI W LOC OF 30 MINUTES OR LESS, SEQUELA
C2832058|T037|S06.301A|ICD10CM|UNSPECIFIED FOCAL TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|UNSP FOCAL TBI W LOC OF 30 MINUTES OR LESS, INIT
C2888900|T047|M00.822|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, LEFT ELBOW|ARTHRITIS DUE TO OTHER BACTERIA, LEFT ELBOW
C2888899|T047|M00.821|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, RIGHT ELBOW|ARTHRITIS DUE TO OTHER BACTERIA, RIGHT ELBOW
C2837743|T037|S32.132A|ICD10CM|SEVERELY DISPLACED ZONE III FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SEVERELY DISPLACED ZONE III FRACTURE OF SACRUM, INIT
C2837744|T037|S32.132B|ICD10CM|SEVERELY DISPLACED ZONE III FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|SEVERELY DISPLACED ZONE III FX SACRUM, INIT FOR OPN FX
C2888901|T047|M00.829|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, UNSPECIFIED ELBOW|ARTHRITIS DUE TO OTHER BACTERIA, UNSPECIFIED ELBOW
C2931826|T047|G71.19|ICD10CM|OTHER SPECIFIED MYOTONIC DISORDERS|MYOTONIA PERMANENS
C2874690|T048|F16.180|ICD10CM|HALLUCINOGEN ABUSE WITH HALLUCINOGEN-INDUCED ANXIETY DISORDER|HALLUCINOGEN ABUSE W HALLUCINOGEN-INDUCED ANXIETY DISORDER
C2874689|T048|F16.188|ICD10CM|HALLUCINOGEN ABUSE WITH OTHER HALLUCINOGEN-INDUCED DISORDER|HALLUCINOGEN ABUSE WITH OTHER HALLUCINOGEN-INDUCED DISORDER
C2885901|T037|T63.832A|ICD10CM|TOXIC EFFECT OF CONTACT WITH OTHER VENOMOUS AMPHIBIAN, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CONTACT W OTH VENOMOUS AMPHIB, SLF-HRM, INIT
C2887768|T047|K50.118|ICD10CM|CROHN'S DISEASE OF LARGE INTESTINE WITH OTHER COMPLICATION|CROHN'S DISEASE OF LARGE INTESTINE WITH OTHER COMPLICATION
C2887769|T047|K50.119|ICD10CM|CROHN'S DISEASE OF LARGE INTESTINE WITH UNSPECIFIED COMPLICATIONS|CROHN'S DISEASE OF LARGE INTESTINE WITH UNSP COMPLICATIONS
C2835212|T037|S22.018B|ICD10CM|OTHER FRACTURE OF FIRST THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF FIRST THORACIC VERTEBRA, INIT FOR OPN FX
C2887767|T047|K50.114|ICD10CM|CROHN'S DISEASE OF LARGE INTESTINE WITH ABSCESS|CROHN'S DISEASE OF LARGE INTESTINE WITH ABSCESS
C2885903|T037|T63.832S|ICD10CM|TOXIC EFFECT OF CONTACT WITH OTHER VENOMOUS AMPHIBIAN, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CONTACT W OTH VENOM AMPHIB, SLF-HRM, SEQUELA
C2887764|T047|K50.111|ICD10CM|CROHN'S DISEASE OF LARGE INTESTINE WITH RECTAL BLEEDING|CROHN'S DISEASE OF LARGE INTESTINE WITH RECTAL BLEEDING
C2887765|T047|K50.112|ICD10CM|CROHN'S DISEASE OF LARGE INTESTINE WITH INTESTINAL OBSTRUCTION|CROHN'S DISEASE OF LARGE INTESTINE W INTESTINAL OBSTRUCTION
C2887766|T047|K50.113|ICD10CM|CROHN'S DISEASE OF LARGE INTESTINE WITH FISTULA|CROHN'S DISEASE OF LARGE INTESTINE WITH FISTULA
C4268182|T047|E66.2|ICD10CM|MORBID (SEVERE) OBESITY WITH ALVEOLAR HYPOVENTILATION|OBESITY HYPOVENTILATION SYNDROME (OHS)
C2858201|T037|S72.365C|ICD10CM|NONDISPLACED SEGMENTAL FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP SEG FX SHAFT OF L FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2858200|T037|S72.365B|ICD10CM|NONDISPLACED SEGMENTAL FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP SEG FX SHAFT OF L FEMUR, INIT FOR OPN FX TYPE I/2
C2858199|T037|S72.365A|ICD10CM|NONDISPLACED SEGMENTAL FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED SEGMENTAL FRACTURE OF SHAFT OF LEFT FEMUR, INIT
C2910916|T033|Z48.22|ICD10CM|ENCOUNTER FOR AFTERCARE FOLLOWING KIDNEY TRANSPLANT|ENCOUNTER FOR AFTERCARE FOLLOWING KIDNEY TRANSPLANT
C2877789|T037|T40.8X2A|ICD10CM|POISONING BY LYSERGIDE [LSD], INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY LYSERGIDE, INTENTIONAL SELF-HARM, INIT ENCNTR
C2888397|T047|L89.221|ICD10CM|PRESSURE ULCER OF LEFT HIP, STAGE 1|PRESSURE ULCER OF LEFT HIP, STAGE 1
C2931689|T047||ICD10CM|MYOTONIC MUSCULAR DYSTROPHY
C2888403|T047|L89.223|ICD10CM|PRESSURE ULCER OF LEFT HIP, STAGE 3|PRESSURE ULCER OF LEFT HIP, STAGE 3
C2888400|T047|L89.222|ICD10CM|PRESSURE ULCER OF LEFT HIP, STAGE 2|PRESSURE ULCER OF LEFT HIP, STAGE 2
C2888406|T047|L89.224|ICD10CM|PRESSURE ULCER OF LEFT HIP, STAGE 4|PRESSURE ULCER OF LEFT HIP, STAGE 4
C2888409|T047|L89.229|ICD10CM|PRESSURE ULCER OF LEFT HIP, UNSPECIFIED STAGE|PRESSURE ULCER OF LEFT HIP, UNSPECIFIED STAGE
C2877791|T037|T40.8X2S|ICD10CM|POISONING BY LYSERGIDE [LSD], INTENTIONAL SELF-HARM, SEQUELA|POISONING BY LYSERGIDE [LSD], INTENTIONAL SELF-HARM, SEQUELA
C2833653|T037|S12.9XXA|ICD10CM|FRACTURE OF NECK, UNSPECIFIED, INITIAL ENCOUNTER|FRACTURE OF NECK, UNSPECIFIED, INITIAL ENCOUNTER
C2901053|T046|M84.469A|ICD10CM|PATHOLOGICAL FRACTURE, UNSPECIFIED TIBIA AND FIBULA, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, UNSP TIBIA AND FIBULA, INIT FOR FX
C2838051|T037|S32.421B|ICD10CM|DISPLACED FRACTURE OF POSTERIOR WALL OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISP FX OF POSTERIOR WALL OF RIGHT ACETAB, INIT FOR OPN FX
C2880077|T037|T48.5X2S|ICD10CM|POISONING BY OTHER ANTI-COMMON-COLD DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH ANTI-COMMON-COLD DRUGS, SELF-HARM, SEQUELA
C2838050|T037|S32.421A|ICD10CM|DISPLACED FRACTURE OF POSTERIOR WALL OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF POSTERIOR WALL OF RIGHT ACETABULUM, INIT
C2838286|T037|S32.474A|ICD10CM|NONDISPLACED FRACTURE OF MEDIAL WALL OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF MEDIAL WALL OF RIGHT ACETABULUM, INIT
C2838287|T037|S32.474B|ICD10CM|NONDISPLACED FRACTURE OF MEDIAL WALL OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP FX OF MEDIAL WALL OF RIGHT ACETAB, INIT FOR OPN FX
C2882475|T047|I69.069|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING UNSPECIFIED SIDE|OTH PARALYTIC SYNDROME FOL NTRM SUBARACH HEMOR AFF UNSP SIDE
C2882473|T047|I69.064|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING LEFT NON-DOMINANT SIDE|OTH PARLYT SYND FOL NTRM SUBARACH HEMOR AFF LEFT NONDOM SIDE
C2882474|T047|I69.065|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE, BILATERAL|OTH PARALYTIC SYNDROME FOLLOWING NTRM SUBARACH HEMOR, BI
C2882471|T047|I69.062|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING LEFT DOMINANT SIDE|OTH PARLYT SYND FOL NTRM SUBARACH HEMOR AFF LEFT DOM SIDE
C2882472|T047|I69.063|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING RIGHT NON-DOMINANT SIDE|OTH PARLYT SYND FOL NTRM SUBARACH HEMOR AFF R NONDOM SIDE
C2880051|T037|T48.4X2S|ICD10CM|POISONING BY EXPECTORANTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY EXPECTORANTS, INTENTIONAL SELF-HARM, SEQUELA
C2882470|T047|I69.061|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING RIGHT DOMINANT SIDE|OTH PARLYT SYND FOL NTRM SUBARACH HEMOR AFF RIGHT DOM SIDE
C2880075|T037|T48.5X2A|ICD10CM|POISONING BY OTHER ANTI-COMMON-COLD DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH ANTI-COMMON-COLD DRUGS, SELF-HARM, INIT
C2845959|T191|C78.02|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF LEFT LUNG|SECONDARY MALIGNANT NEOPLASM OF LEFT LUNG
C2845958|T191|C78.01|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF RIGHT LUNG|SECONDARY MALIGNANT NEOPLASM OF RIGHT LUNG
C2845957|T191|C78.00|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF UNSPECIFIED LUNG|SECONDARY MALIGNANT NEOPLASM OF UNSPECIFIED LUNG
C2880049|T037|T48.4X2A|ICD10CM|POISONING BY EXPECTORANTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY EXPECTORANTS, INTENTIONAL SELF-HARM, INIT
C1332148|T191||ICD10CM|ACUTE ERYTHROID LEUKEMIA, IN REMISSION
C2976785|T191|C94.00|ICD10CM|ACUTE ERYTHROID LEUKEMIA, NOT HAVING ACHIEVED REMISSION|ACUTE ERYTHROID LEUKEMIA WITH FAILED REMISSION
C2890980|T037|T85.128A|ICD10CM|DISPLACEMENT OF OTHER IMPLANTED ELECTRONIC STIMULATOR OF NERVOUS SYSTEM, INITIAL ENCOUNTER|DISPLACMNT OF IMPLNT ELECTRNC STIMULTR OF NERVOUS SYS, INIT
C2861632|T191|C94.02|ICD10CM|ACUTE ERYTHROID LEUKEMIA, IN RELAPSE|ACUTE ERYTHROID LEUKEMIA, IN RELAPSE
C2884562|T037|T56.6X2S|ICD10CM|TOXIC EFFECT OF TIN AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF TIN AND ITS COMPOUNDS, SELF-HARM, SEQUELA
C2859240|T037|S73.042A|ICD10CM|CENTRAL SUBLUXATION OF LEFT HIP, INITIAL ENCOUNTER|CENTRAL SUBLUXATION OF LEFT HIP, INITIAL ENCOUNTER
C2878974|T037|T44.902A|ICD10CM|POISONING BY UNSPECIFIED DRUGS PRIMARILY AFFECTING THE AUTONOMIC NERVOUS SYSTEM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY UNSP DRUGS AFF THE AUTONM NRV SYS, SLF-HRM, INIT
C2842063|T191|C4A.51|ICD10CM|MERKEL CELL CARCINOMA OF ANAL SKIN|MERKEL CELL CARCINOMA OF ANAL SKIN
C2884560|T037|T56.6X2A|ICD10CM|TOXIC EFFECT OF TIN AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF TIN AND ITS COMPOUNDS, SELF-HARM, INIT
C2853900|T191|C83.16|ICD10CM|MANTLE CELL LYMPHOMA, INTRAPELVIC LYMPH NODES|MANTLE CELL LYMPHOMA, INTRAPELVIC LYMPH NODES
C2018777|T191||ICD10CM|MANTLE CELL LYMPHOMA, SPLEEN
C2853898|T191|C83.14|ICD10CM|MANTLE CELL LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB|MANTLE CELL LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB
C2853899|T191|C83.15|ICD10CM|MANTLE CELL LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|MANTLE CELL LYMPHOMA, NODES OF ING REGION AND LOWER LIMB
C2853896|T191|C83.12|ICD10CM|MANTLE CELL LYMPHOMA, INTRATHORACIC LYMPH NODES|MANTLE CELL LYMPHOMA, INTRATHORACIC LYMPH NODES
C2853897|T191|C83.13|ICD10CM|MANTLE CELL LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES|MANTLE CELL LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES
C2873962|T047|E09.29|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH OTHER DIABETIC KIDNEY COMPLICATION|DRUG/CHEM DIABETES W OTH DIABETIC KIDNEY COMPLICATION
C2853895|T191|C83.11|ICD10CM|MANTLE CELL LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK|MANTLE CELL LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK
C2873960|T047|E09.22|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH DIABETIC CHRONIC KIDNEY DISEASE|DRUG/CHEM DIABETES W DIABETIC CHRONIC KIDNEY DISEASE
C2873959|T047|E09.21|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH DIABETIC NEPHROPATHY|DRUG/CHEM DIABETES MELLITUS W DIABETIC NEPHROPATHY
C2887937|T047|K72.91|ICD10CM|HEPATIC FAILURE, UNSPECIFIED WITH COMA|HEPATIC FAILURE, UNSPECIFIED WITH COMA
C2848460|T037|S58.922S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT FOREARM, LEVEL UNSPECIFIED, SEQUELA|PARTIAL TRAUMATIC AMP OF L FOREARM, LEVEL UNSP, SEQUELA
C2889919|T037|T82.321A|ICD10CM|DISPLACEMENT OF CAROTID ARTERIAL GRAFT (BYPASS), INITIAL ENCOUNTER|DISPLACEMENT OF CAROTID ARTERIAL GRAFT (BYPASS), INIT ENCNTR
C2833323|T037|S12.201A|ICD10CM|UNSPECIFIED NONDISPLACED FRACTURE OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP NONDISP FX OF THIRD CERVICAL VERTEBRA, INIT FOR CLOS FX
C2833324|T037|S12.201B|ICD10CM|UNSPECIFIED NONDISPLACED FRACTURE OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP NONDISP FX OF THIRD CERVICAL VERTEBRA, INIT FOR OPN FX
C2834013|T037|S14.146A|ICD10CM|BROWN-SEQUARD SYNDROME AT C6 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|BROWN-SEQUARD SYNDROME AT C6, INIT
C0260764|T033|Z43.4|DMDICD10|ENCOUNTER FOR ATTENTION TO OTHER ARTIFICIAL OPENINGS OF DIGESTIVE TRACT|VERSORGUNG ANDERER KUENSTLICHER KOERPEROEFFNUNGEN DES VERDAUUNGSTRAKTES
C4269496|T037|S02.632A|ICD10CM|FRACTURE OF CORONOID PROCESS OF LEFT MANDIBLE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF CORONOID PROCESS OF LEFT MANDIBLE, INIT
C2901147|T046|M84.512A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, LEFT SHOULDER, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, L SHOULDER, INIT
C2901871|T047|M86.421|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, RIGHT HUMERUS|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, RIGHT HUMERUS
C2901872|T047|M86.422|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, LEFT HUMERUS|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, LEFT HUMERUS
C2901873|T047|M86.429|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, UNSPECIFIED HUMERUS|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, UNSP HUMERUS
C0740203|T033|Z43|DMDICD10|ENCOUNTER FOR ATTENTION TO UNSPECIFIED ARTIFICIAL OPENING|VERSORGUNG KUENSTLICHER KOERPEROEFFNUNGEN
C4269501|T037|S02.632S|ICD10CM|FRACTURE OF CORONOID PROCESS OF LEFT MANDIBLE, SEQUELA|FRACTURE OF CORONOID PROCESS OF LEFT MANDIBLE, SEQUELA
C4268260|T048|F15.988|ICD10CM|OTHER STIMULANT USE, UNSPECIFIED WITH OTHER STIMULANT-INDUCED DISORDER|AMPHETAMINE OR OTHER STIMULANT-INDUCED OBSESSIVE COMPULSIVE OR RELATED DISORDER, WITHOUT USE DISORDER
C2832559|T037|S06.812S|ICD10CM|INJURY OF RIGHT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|INJURY OF R INT CAROTID, INTCR W LOC OF 31-59 MIN, SEQUELA
C4237016|T048|F15.982|ICD10CM|OTHER STIMULANT USE, UNSPECIFIED WITH STIMULANT-INDUCED SLEEP DISORDER|CAFFEINE INDUCED SLEEP DISORDER, WITHOUT USE DISORDER
C4236977|T048|F15.981|ICD10CM|OTHER STIMULANT USE, UNSPECIFIED WITH STIMULANT-INDUCED SEXUAL DYSFUNCTION|AMPHETAMINE OR OTHER STIMULANT-INDUCED SEXUAL DYSFUNCTION, WITHOUT USE DISORDER
C0348362|T191|C49.9|DMDICD10|MALIGNANT NEOPLASM OF CONNECTIVE AND SOFT TISSUE, UNSPECIFIED|BOESARTIGE NEUBILDUNG: BINDEGEWEBE UND ANDERE WEICHTEILGEWEBE, NICHT NAEHER BEZEICHNET
C2874588|T048|F14.19|ICD10CM|COCAINE ABUSE WITH UNSPECIFIED COCAINE-INDUCED DISORDER|COCAINE ABUSE WITH UNSPECIFIED COCAINE-INDUCED DISORDER
C2901401|T046|M84.622A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, LEFT HUMERUS, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, LEFT HUMERUS, INIT
C2832465|T037|S06.4X9A|ICD10CM|EPIDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|EPIDURAL HEMORRHAGE W LOC OF UNSP DURATION, INIT
C2865559|T037|S88.122A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, LEFT LOWER LEG, INITIAL ENCOUNTER|PART TRAUM AMP AT LEVEL BETW KNEE AND ANKLE, L LOW LEG, INIT
C2874513|T048|F13.120|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE WITH INTOXICATION, UNCOMPLICATED|SEDATV/HYP/ANXIOLYTC ABUSE W INTOXICATION, UNCOMPLICATED
C2865560|T037|S88.122D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, LEFT LOWER LEG, SUBSEQUENT ENCOUNTER|PART TRAUM AMP AT LEVEL BETW KNEE AND ANKLE, L LOW LEG, SUBS
C2888825|T047||ICD10CM|STAPHYLOCOCCAL ARTHRITIS, VERTEBRAE
C2888826|T047|M00.09|ICD10CM|STAPHYLOCOCCAL POLYARTHRITIS|STAPHYLOCOCCAL POLYARTHRITIS
C0260686|T033|Z93.4|DMDICD10|OTHER ARTIFICIAL OPENINGS OF GASTROINTESTINAL TRACT STATUS|VORHANDENSEIN ANDERER KUENSTLICHER KOERPEROEFFNUNGEN DES MAGEN-DARMTRAKTES
C0260684|T033|Z93.2|DMDICD10|ILEOSTOMY STATUS|VORHANDENSEIN EINES ILEOSTOMAS
C0260685|T033|Z93.3|DMDICD10|COLOSTOMY STATUS|VORHANDENSEIN EINES KOLOSTOMAS
C0260682|T033|Z93.0|DMDICD10|TRACHEOSTOMY STATUS|VORHANDENSEIN EINES TRACHEOSTOMAS
C0260683|T033|Z93.1|DMDICD10|GASTROSTOMY STATUS|VORHANDENSEIN EINES GASTROSTOMAS
C2888793|T047|M00.00|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, UNSPECIFIED JOINT|STAPHYLOCOCCAL ARTHRITIS, UNSPECIFIED JOINT
C2832467|T037|S06.4X9S|ICD10CM|EPIDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|EPIDURAL HEMORRHAGE W LOC OF UNSP DURATION, SEQUELA
C2857139|T037|S72.109C|ICD10CM|UNSPECIFIED TROCHANTERIC FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP TROCHAN FX UNSP FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2857138|T037|S72.109B|ICD10CM|UNSPECIFIED TROCHANTERIC FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP TROCHAN FX UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2857137|T037|S72.109A|ICD10CM|UNSPECIFIED TROCHANTERIC FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP TROCHANTERIC FRACTURE OF UNSP FEMUR, INIT FOR CLOS FX
C0260691|T033|Z93|DMDICD10|ARTIFICIAL OPENING STATUS, UNSPECIFIED|VORHANDENSEIN EINER KUENSTLICHEN KOERPEROEFFNUNG
C2889562|T047|M08.242|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, LEFT HAND|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, LEFT HAND
C2889561|T047|M08.241|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, RIGHT HAND|JUVENILE RHEUMATOID ARTHRITIS W SYSTEMIC ONSET, RIGHT HAND
C2884416|T037|T54.92XS|ICD10CM|TOXIC EFFECT OF UNSPECIFIED CORROSIVE SUBSTANCE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF UNSP CORROSIVE SUBSTANCE, SELF-HARM, SEQUELA
C2889560|T047|M08.24|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, UNSPECIFIED HAND|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, HAND
C2874765|T048|F18.250|ICD10CM|INHALANT DEPENDENCE WITH INHALANT-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|INHALANT DEPEND W INHALNT-INDUCE PSYCH DISORDER W DELUSIONS
C2874766|T048|F18.251|ICD10CM|INHALANT DEPENDENCE WITH INHALANT-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|INHALANT DEPEND W INHALNT-INDUCE PSYCH DISORDER W HALLUCIN
C2874767|T048|F18.259|ICD10CM|INHALANT DEPENDENCE WITH INHALANT-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|INHALANT DEPENDENCE WITH INHALANT-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED
C2888867|T047|M00.229|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, UNSPECIFIED ELBOW|OTHER STREPTOCOCCAL ARTHRITIS, UNSPECIFIED ELBOW
C2888865|T047|M00.221|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, RIGHT ELBOW|OTHER STREPTOCOCCAL ARTHRITIS, RIGHT ELBOW
C2888866|T047|M00.222|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, LEFT ELBOW|OTHER STREPTOCOCCAL ARTHRITIS, LEFT ELBOW
C0348988|T047|B52.0|DMDICD10|PLASMODIUM MALARIAE MALARIA WITH NEPHROPATHY|MALARIA QUARTANA MIT NEPHROPATHIE
C2889530|T047|M08.022|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, LEFT ELBOW|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, LEFT ELBOW
C2889529|T047|M08.021|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, RIGHT ELBOW|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, RIGHT ELBOW
C2832561|T037|S06.813A|ICD10CM|INJURY OF RIGHT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|INJURY OF R INT CAROTID, INTCR W LOC OF 1-5 HRS 59 MIN, INIT
C2889531|T047|M08.02|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED ELBOW|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS OF ELBOW
C2876743|T037|T36.8X2A|ICD10CM|POISONING BY OTHER SYSTEMIC ANTIBIOTICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH SYSTEMIC ANTIBIOTICS, SELF-HARM, INIT
C4270153|T046|T82.848A|ICD10CM|PAIN DUE TO VASCULAR PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|PAIN DUE TO VASCULAR PROSTH DEV/GRFT, INITIAL ENCOUNTER
C2882370|T047|I63.329|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF UNSPECIFIED ANTERIOR CEREBRAL ARTERY|CEREBRAL INFRC DUE TO THOMBOS UNSP ANTERIOR CEREBRAL ARTERY
C0155918|T047|J98.3|DMDICD10|COMPENSATORY EMPHYSEMA|KOMPENSATORISCHES EMPHYSEM
C1370824|T047|J98.2|DMDICD10|INTERSTITIAL EMPHYSEMA|INTERSTITIELLES EMPHYSEM
C2876149|T037|T31.61|ICD10CM|BURNS INVOLVING 60-69% OF BODY SURFACE WITH 10-19% THIRD DEGREE BURNS|BURNS OF 60-69% OF BODY SURFACE W 10-19% THIRD DEGREE BURNS
C2873891|T047|E08.21|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH DIABETIC NEPHROPATHY|DIABETES DUE TO UNDERLYING CONDITION W DIABETIC NEPHROPATHY
C2876154|T037|T31.66|ICD10CM|BURNS INVOLVING 60-69% OF BODY SURFACE WITH 60-69% THIRD DEGREE BURNS|BURNS OF 60-69% OF BODY SURFACE W 60-69% THIRD DEGREE BURNS
C2876153|T037|T31.65|ICD10CM|BURNS INVOLVING 60-69% OF BODY SURFACE WITH 50-59% THIRD DEGREE BURNS|BURNS OF 60-69% OF BODY SURFACE W 50-59% THIRD DEGREE BURNS
C2876152|T037|T31.64|ICD10CM|BURNS INVOLVING 60-69% OF BODY SURFACE WITH 40-49% THIRD DEGREE BURNS|BURNS OF 60-69% OF BODY SURFACE W 40-49% THIRD DEGREE BURNS
C2878637|T037|T43.632S|ICD10CM|POISONING BY METHYLPHENIDATE, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY METHYLPHENIDATE, INTENTIONAL SELF-HARM, SEQUELA
C2905672|T037|X72.XXXA|ICD10CM|INTENTIONAL SELF-HARM BY HANDGUN DISCHARGE, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY HANDGUN DISCHARGE, INIT ENCNTR
C1561636|T047||ICD10CM|SCLEROSING MESENTERITIS
C2887906|T047|K65.0|ICD10CM|GENERALIZED (ACUTE) PERITONITIS|SUBPHRENIC PERITONITIS (ACUTE)
C0267762|T047|K65.1|ICD10CM|PERITONEAL ABSCESS|SUBHEPATIC ABSCESS
C0275551|T047|K65.2|ICD10CM|SPONTANEOUS BACTERIAL PERITONITIS|SPONTANEOUS BACTERIAL PERITONITIS
C0267768|T047|K65.3|ICD10CM|CHOLEPERITONITIS|PERITONITIS DUE TO BILE
C2842065|T191|C4A.59|ICD10CM|MERKEL CELL CARCINOMA OF OTHER PART OF TRUNK|MERKEL CELL CARCINOMA OF OTHER PART OF TRUNK
C0348746|T047|K65.8|DMDICD10|OTHER PERITONITIS|SONSTIGE PERITONITIS
C0275550|T047||ICD10CM|PERITONITIS, UNSPECIFIED
C0152234|T019|Q00.2|DMDICD10|INIENCEPHALY|INIENZEPHALIE
C4268482|T047|I63.323|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF BILATERAL ANTERIOR CEREBRAL ARTERIES|CEREBRAL INFRC DUE TO THOMBOS OF BI ANT CEREBRAL ARTERIES
C2843321|T037|S48.911A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT SHOULDER AND UPPER ARM, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|COMPLETE TRAUM AMP OF RIGHT SHLDR/UP ARM, LEVEL UNSP, INIT
C2882677|T046|I69.962|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING LEFT DOMINANT SIDE|OTH PARLYT SYND FOL UNSP CEREBVASC DISEASE AFF LEFT DOM SIDE
C2858063|T037|S72.353B|ICD10CM|DISPLACED COMMINUTED FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL COMMNT FX SHAFT OF UNSP FEMR, INIT FOR OPN FX TYPE I/2
C2858064|T037|S72.353C|ICD10CM|DISPLACED COMMINUTED FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL COMMNT FX SHAFT OF UNSP FEMR, 7THC
C2858062|T037|S72.353A|ICD10CM|DISPLACED COMMINUTED FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED COMMINUTED FRACTURE OF SHAFT OF UNSP FEMUR, INIT
C2882368|T047|I63.321|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF RIGHT ANTERIOR CEREBRAL ARTERY|CEREBRAL INFRC DUE TO THOMBOS OF RIGHT ANT CEREBRAL ARTERY
C2831448|T037|S02.119S|ICD10CM|UNSPECIFIED FRACTURE OF OCCIPUT, SEQUELA|UNSPECIFIED FRACTURE OF OCCIPUT, SEQUELA
C0694506|T047|K23|DMDICD10|DISORDERS OF ESOPHAGUS IN DISEASES CLASSIFIED ELSEWHERE|KRANKHEITEN DES OESOPHAGUS BEI ANDERENORTS KLASSIFIZIERTEN KRANKHEITEN
C2855957|T037|S68.419S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED HAND AT WRIST LEVEL, SEQUELA|COMPLETE TRAUMATIC AMP OF UNSP HAND AT WRIST LEVEL, SEQUELA
C2831444|T037|S02.119B|ICD10CM|UNSPECIFIED FRACTURE OF OCCIPUT, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF OCCIPUT, INIT ENCNTR FOR OPEN FRACTURE
C2831443|T037|S02.119A|ICD10CM|UNSPECIFIED FRACTURE OF OCCIPUT, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF OCCIPUT, INIT ENCNTR FOR CLOSED FRACTURE
C2869843|T037|S98.219D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF TWO OR MORE UNSPECIFIED LESSER TOES, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMP OF TWO OR MORE UNSP LESSER TOES, SUBS
C2855955|T037|S68.419A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED HAND AT WRIST LEVEL, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMP OF UNSP HAND AT WRIST LEVEL, INIT
C0154050|T191||ICD10AM|HEMANGIOMA OF INTRACRANIAL STRUCTURES
C2901986|T046|M87.111|ICD10CM|OSTEONECROSIS DUE TO DRUGS, RIGHT SHOULDER|OSTEONECROSIS DUE TO DRUGS, RIGHT SHOULDER
C0003873|T047|M06.9|DMDICD10|RHEUMATOID ARTHRITIS, UNSPECIFIED|CHRONISCHE POLYARTHRITIS, NICHT NAEHER BEZEICHNET
C2874792|T048|F19.120|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE ABUSE WITH INTOXICATION, UNCOMPLICATED|OTH PSYCHOACTIVE SUBSTANCE ABUSE W INTOXICATION, UNCOMP
C2874794|T048|F19.122|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE ABUSE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCES|OTH PSYCHOACTV SUBSTANCE ABUSE W INTOX W PERCEPTUAL DISTURB
C0162323|T047|M13.0|DMDICD10|INFLAMMATORY POLYARTHROPATHY|POLYARTHRITIS, NICHT NAEHER BEZEICHNET
C2901502|T046|M84.659A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, HIP, UNSPECIFIED, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, HIP, UNSP, INIT FOR FX
C2874795|T048|F19.12|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE ABUSE WITH INTOXICATION, UNSPECIFIED|OTHER PSYCHOACTIVE SUBSTANCE ABUSE WITH INTOXICATION
C0839946|T047|M86.18|ICD10AM|OTHER ACUTE OSTEOMYELITIS, OTHER SITE|OTHER ACUTE OSTEOMYELITIS, OTHER SITE
C3263903|T037|T81.12XA|ICD10CM|POSTPROCEDURAL SEPTIC SHOCK, INITIAL ENCOUNTER|POSTPROCEDURAL SEPTIC SHOCK, INITIAL ENCOUNTER
C0343052|T047|L40.4|DMDICD10|GUTTATE PSORIASIS|PSORIASIS GUTTATA
C2885341|T037|T63.022S|ICD10CM|TOXIC EFFECT OF CORAL SNAKE VENOM, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CORAL SNAKE VENOM, SELF-HARM, SEQUELA
C0406317|T047|L40.0|ICD10CM|PSORIASIS VULGARIS|NUMMULAR PSORIASIS
C2888177|T047|L40.1|ICD10CM|GENERALIZED PUSTULAR PSORIASIS|VON ZUMBUSCH'S DISEASE
C0392439|T047|L40.2|DMDICD10|ACRODERMATITIS CONTINUA|AKRODERMATITIS CONTINUA SUPPURATIVA [HALLOPEAU]
C0030246|T047|L40.3|DMDICD10|PUSTULOSIS PALMARIS ET PLANTARIS|PSORIASIS PUSTULOSA PALMOPLANTARIS
C0477485|T047|L40.8|DMDICD10|OTHER PSORIASIS|SONSTIGE PSORIASIS
C0033860|T047|L40.9|DMDICD10|PSORIASIS, UNSPECIFIED|PSORIASIS, NICHT NAEHER BEZEICHNET
C0267088|T020||ICD10CM|DIVERTICULUM OF ESOPHAGUS, ACQUIRED
C2889094|T047|M02.851|ICD10CM|OTHER REACTIVE ARTHROPATHIES, RIGHT HIP|OTHER REACTIVE ARTHROPATHIES, RIGHT HIP
C2889095|T047|M02.852|ICD10CM|OTHER REACTIVE ARTHROPATHIES, LEFT HIP|OTHER REACTIVE ARTHROPATHIES, LEFT HIP
C1321756|T047||ICD10CM|ACHALASIA OF CARDIA
C0281839|T037|K22.3|ICD10CM|PERFORATION OF ESOPHAGUS|RUPTURE OF ESOPHAGUS
C1393788|T020||ICD10CM|ESOPHAGEAL OBSTRUCTION
C2362829|T191|C48.1|ICD10CM|MALIGNANT NEOPLASM OF SPECIFIED PARTS OF PERITONEUM|MALIGNANT NEOPLASM OF PELVIC PERITONEUM
C2889096|T047|M02.85|ICD10CM|OTHER REACTIVE ARTHROPATHIES, UNSPECIFIED HIP|OTHER REACTIVE ARTHROPATHIES, HIP
C2858695|T037|S72.444A|ICD10CM|NONDISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF LOWER EPIPHYSIS (SEPARATION) OF R FEMUR, INIT
C0153467|T191|C48.2|DMDICD10|MALIGNANT NEOPLASM OF PERITONEUM, UNSPECIFIED|BOESARTIGE NEUBILDUNG: PERITONEUM, NICHT NAEHER BEZEICHNET
C0014852|T047|K22.9|DMDICD10|DISEASE OF ESOPHAGUS, UNSPECIFIED|KRANKHEIT DES OESOPHAGUS, NICHT NAEHER BEZEICHNET
C0348727|T047|K22.8|DMDICD10|OTHER SPECIFIED DISEASES OF ESOPHAGUS|SONSTIGE NAEHER BEZEICHNETE KRANKHEITEN DES OESOPHAGUS
C2857086|T037|S72.099B|ICD10CM|OTHER FRACTURE OF HEAD AND NECK OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|OTH FX HEAD/NECK OF UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2882406|T046|I63.529|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF UNSPECIFIED ANTERIOR CEREBRAL ARTERY|CEREB INFRC D/T UNSP OCCLS OR STENOS OF UNSP ANT CEREB ART
C2882404|T046|I63.521|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF RIGHT ANTERIOR CEREBRAL ARTERY|CEREB INFRC D/T UNSP OCCLS OR STENOS OF RIGHT ANT CEREB ART
C4268490|T046|I63.523|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF BILATERAL ANTERIOR CEREBRAL ARTERIES|CEREB INFRC DUE TO UNSP OCCLS OR STENOS OF BI ANT CEREB ART
C2882405|T046|I63.522|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF LEFT ANTERIOR CEREBRAL ARTERY|CEREB INFRC D/T UNSP OCCLS OR STENOS OF LEFT ANT CEREB ART
C2856015|T037|S68.613S|ICD10CM|COMPLETE TRAUMATIC TRANSPHALANGEAL AMPUTATION OF LEFT MIDDLE FINGER, SEQUELA|COMPLETE TRAUMATIC TRNSPHAL AMP OF L MID FINGER, SEQUELA
C4316812|T047||ICD10CM|HEREDITARY DEFICIENCY OF OTHER CLOTTING FACTORS
C4269475|T037|S02.622A|ICD10CM|FRACTURE OF SUBCONDYLAR PROCESS OF LEFT MANDIBLE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF SUBCONDYLAR PROCESS OF LEFT MANDIBLE, INIT
C2845946|T191|C74.90|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED PART OF UNSPECIFIED ADRENAL GLAND|MALIGNANT NEOPLASM OF UNSP PART OF UNSPECIFIED ADRENAL GLAND
C2845947|T191|C74.91|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED PART OF RIGHT ADRENAL GLAND|MALIGNANT NEOPLASM OF UNSP PART OF RIGHT ADRENAL GLAND
C2845948|T191|C74.92|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED PART OF LEFT ADRENAL GLAND|MALIGNANT NEOPLASM OF UNSPECIFIED PART OF LEFT ADRENAL GLAND
C2890642|T037|T84.126A|ICD10CM|DISPLACEMENT OF INTERNAL FIXATION DEVICE OF BONE OF RIGHT LOWER LEG, INITIAL ENCOUNTER|DISPLACEMENT OF INT FIX OF BONE OF RIGHT LOWER LEG, INIT
C3263948|T046|D68.32|ICD10CM|HEMORRHAGIC DISORDER DUE TO EXTRINSIC CIRCULATING ANTICOAGULANTS|HEMORRHAGIC DISORDER DUE TO INCREASE IN ANTI-XA
C2830383|T033|R40.2223|ICD10CM|COMA SCALE, BEST VERBAL RESPONSE, INCOMPREHENSIBLE WORDS, AT HOSPITAL ADMISSION|COMA SCALE, BEST VERB, INCOMPREHENSIBLE WORDS, ADMIT
C2830382|T033|R40.2222|ICD10CM|COMA SCALE, BEST VERBAL RESPONSE, INCOMPREHENSIBLE WORDS, AT ARRIVAL TO EMERGENCY DEPARTMENT|COMA SCALE, BEST VERB, INCOMPREHENSIBLE WORDS, EMR
C2830381|T033|R40.2221|ICD10CM|COMA SCALE, BEST VERBAL RESPONSE, INCOMPREHENSIBLE WORDS, IN THE FIELD [EMT OR AMBULANCE]|COMA SCALE, BEST VERB, INCOMPREHENSIBLE WORDS, IN THE FIELD
C2830380|T033|R40.2220|ICD10CM|COMA SCALE, BEST VERBAL RESPONSE, INCOMPREHENSIBLE WORDS, UNSPECIFIED TIME|COMA SCALE, BEST VERB, INCOMPREHENSIBLE WORDS, UNSP TIME
C2832154|T037|S06.324S|ICD10CM|CONTUSION AND LACERATION OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|CONTUS/LAC LEFT CEREBRUM W LOC OF 6-24 HRS, SEQUELA
C2830384|T033|R40.2224|ICD10CM|COMA SCALE, BEST VERBAL RESPONSE, INCOMPREHENSIBLE WORDS, 24 HOURS OR MORE AFTER HOSPITAL ADMISSION|COMA SCALE, BEST VERB, INCOMPREHENSIBLE WORDS, 24+HRS
C4267989|T047|E09.3532|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, LEFT EYE|DRUG/CHEM DIAB W PROLIF DIAB RTNOP W TRCTN DTCH N-MCLA,L EYE
C4267990|T047|E09.3533|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, BILATERAL|DRUG/CHEM DIAB W PROLIF DIAB RTNOP W TRCTN DTCH N-MCLA, BI
C4267988|T047|E09.3531|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, RIGHT EYE|DRUG/CHEM DIAB W PROLIF DIAB RTNOP W TRCTN DTCH N-MCLA,R EYE
C2832152|T037|S06.324A|ICD10CM|CONTUSION AND LACERATION OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|CONTUS/LAC LEFT CEREBRUM W LOC OF 6 HOURS TO 24 HOURS, INIT
C4267991|T047|E09.3539|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, UNSPECIFIED EYE|DRUG/CHEM DIAB W PROLIF DIAB RTNOP W TRCTN DTCH N-MCLA, UNSP
C2910348|T047||ICD10CM|MARFAN'S SYNDROME WITH SKELETAL MANIFESTATION
C2882874|T047|I70.523|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, BILATERAL LEGS|ATHSCL NONAUT BIO BYPASS OF THE EXTRM W REST PAIN, BI LEGS
C0024796|T047|Q87.40|ICD10CM|MARFAN'S SYNDROME, UNSPECIFIED|MARFAN'S SYNDROME, UNSPECIFIED
C2905807|T037|X83.0XXD|ICD10CM|INTENTIONAL SELF-HARM BY CRASHING OF AIRCRAFT, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY CRASHING OF AIRCRAFT, SUBS ENCNTR
C2879872|T037|T47.8X2S|ICD10CM|POISONING BY OTHER AGENTS PRIMARILY AFFECTING GASTROINTESTINAL SYSTEM, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH AGENTS AFF GI SYS, SELF-HARM, SEQUELA
C2905806|T037|X83.0XXA|ICD10CM|INTENTIONAL SELF-HARM BY CRASHING OF AIRCRAFT, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY CRASHING OF AIRCRAFT, INIT ENCNTR
C2832012|T037|S06.2X0A|ICD10CM|DIFFUSE TRAUMATIC BRAIN INJURY WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|DIFFUSE TBI W/O LOSS OF CONSCIOUSNESS, INIT
C0011302|T047|G37.9|DMDICD10|DEMYELINATING DISEASE OF CENTRAL NERVOUS SYSTEM, UNSPECIFIED|DEMYELINISIERENDE KRANKHEIT DES ZENTRALNERVENSYSTEMS, NICHT NAEHER BEZEICHNET
C0393663|T047|G37.8|DMDICD10|OTHER SPECIFIED DEMYELINATING DISEASES OF CENTRAL NERVOUS SYSTEM|SONSTIGE NAEHER BEZEICHNETE DEMYELINISIERENDE KRANKHEITEN DES ZENTRALNERVENSYSTEMS
C2905808|T037|X83.0XXS|ICD10CM|INTENTIONAL SELF-HARM BY CRASHING OF AIRCRAFT, SEQUELA|INTENTIONAL SELF-HARM BY CRASHING OF AIRCRAFT, SEQUELA
C2875071|T047|G37.3|ICD10CM|ACUTE TRANSVERSE MYELITIS IN DEMYELINATING DISEASE OF CENTRAL NERVOUS SYSTEM|ACUTE TRANSVERSE MYELOPATHY
C0206083|T047|G37.2|DMDICD10|CENTRAL PONTINE MYELINOLYSIS|ZENTRALE PONTINE MYELINOLYSE
C0238265|T047|G37.1|DMDICD10|CENTRAL DEMYELINATION OF CORPUS CALLOSUM|ZENTRALE DEMYELINISATION DES CORPUS CALLOSUM
C2875070|T047||ICD10CM|DIFFUSE SCLEROSIS OF CENTRAL NERVOUS SYSTEM
C2875073|T047|G37.5|ICD10CM|CONCENTRIC SCLEROSIS [BALO] OF CENTRAL NERVOUS SYSTEM|CONCENTRIC SCLEROSIS [BALO] OF CENTRAL NERVOUS SYSTEM
C2875072|T047|G37.4|ICD10CM|SUBACUTE NECROTIZING MYELITIS OF CENTRAL NERVOUS SYSTEM|SUBACUTE NECROTIZING MYELITIS OF CENTRAL NERVOUS SYSTEM
C2895194|T047|M33.99|ICD10CM|DERMATOPOLYMYOSITIS, UNSPECIFIED WITH OTHER ORGAN INVOLVEMENT|DERMATOPOLYMYOSITIS, UNSP WITH OTHER ORGAN INVOLVEMENT
C0236830|T047||ICD10CM|NEUROLEPTIC INDUCED PARKINSONISM
C2882179|T047|I25.710|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN CORONARY ARTERY BYPASS GRAFT(S) WITH UNSTABLE ANGINA PECTORIS|ATHSCL AUTOLOGOUS VEIN CABG W UNSTABLE ANGINA PECTORIS
C2882180|T047|I25.711|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN CORONARY ARTERY BYPASS GRAFT(S) WITH ANGINA PECTORIS WITH DOCUMENTED SPASM|ATHSCL AUTOLOGOUS VEIN CABG W ANG PCTRS W DOCUMENTED SPASM
C2895192|T047|M33.91|ICD10CM|DERMATOPOLYMYOSITIS, UNSPECIFIED WITH RESPIRATORY INVOLVEMENT|DERMATOPOLYMYOSITIS, UNSP WITH RESPIRATORY INVOLVEMENT
C0011633|T047|M33.90|ICD10CM|DERMATOPOLYMYOSITIS, UNSPECIFIED, ORGAN INVOLVEMENT UNSPECIFIED|DERMATOPOLYMYOSITIS, UNSPECIFIED, ORGAN INVOLVEMENT UNSPECIFIED
C4509354|T047|M33.93|ICD10CM|DERMATOPOLYMYOSITIS, UNSPECIFIED WITHOUT MYOPATHY|DERMATOPOLYMYOSITIS, UNSPECIFIED WITHOUT MYOPATHY
C4237315|T047|G21.19|ICD10CM|OTHER DRUG INDUCED SECONDARY PARKINSONISM|OTHER MEDICATION-INDUCED PARKINSONISM
C2882181|T047|I25.718|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN CORONARY ARTERY BYPASS GRAFT(S) WITH OTHER FORMS OF ANGINA PECTORIS|ATHSCL AUTOLOGOUS VEIN CABG W OTH ANGINA PECTORIS
C2882182|T047|I25.719|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN CORONARY ARTERY BYPASS GRAFT(S) WITH UNSPECIFIED ANGINA PECTORIS|ATHSCL AUTOLOGOUS VEIN CABG W UNSP ANGINA PECTORIS
C2890414|T037|T84.013A|ICD10CM|BROKEN INTERNAL LEFT KNEE PROSTHESIS, INITIAL ENCOUNTER|BROKEN INTERNAL LEFT KNEE PROSTHESIS, INITIAL ENCOUNTER
C2838351|T037|S32.491A|ICD10CM|OTHER SPECIFIED FRACTURE OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF RIGHT ACETABULUM, INIT FOR CLOS FX
C2837999|T191|C43.62|ICD10CM|MALIGNANT MELANOMA OF LEFT UPPER LIMB, INCLUDING SHOULDER|MALIGNANT MELANOMA OF LEFT UPPER LIMB, INCLUDING SHOULDER
C2837998|T191|C43.61|ICD10CM|MALIGNANT MELANOMA OF RIGHT UPPER LIMB, INCLUDING SHOULDER|MALIGNANT MELANOMA OF RIGHT UPPER LIMB, INCLUDING SHOULDER
C2837997|T191|C43.60|ICD10CM|MALIGNANT MELANOMA OF UNSPECIFIED UPPER LIMB, INCLUDING SHOULDER|MALIGNANT MELANOMA OF UNSP UPPER LIMB, INCLUDING SHOULDER
C2886962|T037|T81.522S|ICD10CM|OBSTRUCTION DUE TO FOREIGN BODY ACCIDENTALLY LEFT IN BODY FOLLOWING KIDNEY DIALYSIS, SEQUELA|OBST DUE TO FB ACC LEFT IN BODY FOL KIDNEY DIALYSIS, SEQUELA
C4267921|T047|E08.3511|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|DIAB WITH PROLIF DIABETIC RTNOP WITH MACULAR EDEMA, R EYE
C4267923|T047|E08.3513|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|DIABETES WITH PROLIF DIABETIC RTNOP WITH MACULAR EDEMA, BI
C4267922|T047|E08.3512|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|DIAB WITH PROLIF DIABETIC RTNOP WITH MACULAR EDEMA, LEFT EYE
C4270443|T046|T83.85XA|ICD10CM|STENOSIS DUE TO GENITOURINARY PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|STENOSIS DUE TO GENITOURINARY PROSTH DEV/GRFT, INIT
C4267924|T047|E08.3519|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|DIABETES WITH PROLIF DIABETIC RTNOP WITH MACULAR EDEMA, UNSP
C2837518|T037|S32.020B|ICD10CM|WEDGE COMPRESSION FRACTURE OF SECOND LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|WEDGE COMPRSN FX SECOND LUM VERTEBRA, INIT FOR OPN FX
C2853957|T191|C84.19|ICD10CM|SEZARY DISEASE, EXTRANODAL AND SOLID ORGAN SITES|SÉZARY DISEASE, EXTRANODAL AND SOLID ORGAN SITES
C0153817|T191||ICD10CM|SEZARY DISEASE, LYMPH NODES OF MULTIPLE SITES
C0153810|T191||ICD10CM|SEZARY DISEASE, LYMPH NODES OF HEAD, FACE, AND NECK
C0036920|T191|C84.10|ICD10CM|SEZARY DISEASE, UNSPECIFIED SITE|SÉZARY DISEASE, UNSPECIFIED SITE
C0153812|T191||ICD10CM|SEZARY DISEASE, INTRA-ABDOMINAL LYMPH NODES
C0153811|T191||ICD10CM|SEZARY DISEASE, INTRATHORACIC LYMPH NODES
C0153814|T191|C84.15|ICD10CM|SEZARY DISEASE, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|SEZARY DISEASE, NODES OF INGUINAL REGION AND LOWER LIMB
C0153813|T191||ICD10CM|SEZARY DISEASE, LYMPH NODES OF AXILLA AND UPPER LIMB
C0153816|T191||ICD10CM|SEZARY DISEASE, SPLEEN
C0153815|T191||ICD10CM|SEZARY DISEASE, INTRAPELVIC LYMPH NODES
C4269536|T037|S02.651S|ICD10CM|FRACTURE OF ANGLE OF RIGHT MANDIBLE, SEQUELA|FRACTURE OF ANGLE OF RIGHT MANDIBLE, SEQUELA
C2832393|T037|S06.381S|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF BRAINSTEM WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|CONTUS/LAC/HEM BRNST W LOC OF 30 MINUTES OR LESS, SEQUELA
C2888806|T047|M00.039|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, UNSPECIFIED WRIST|STAPHYLOCOCCAL ARTHRITIS, UNSPECIFIED WRIST
C2349281|T191||ICD10CM|MYELOID SARCOMA, IN RELAPSE
C2861590|T191||ICD10CM|MYELOID SARCOMA, NOT HAVING ACHIEVED REMISSION
C0153892|T191|C92.31|ICD10AM|MYELOID SARCOMA, IN REMISSION|MYELOID SARCOMA, IN REMISSION, IN REMISSION
C2888804|T047|M00.031|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, RIGHT WRIST|STAPHYLOCOCCAL ARTHRITIS, RIGHT WRIST
C2888805|T047|M00.032|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, LEFT WRIST|STAPHYLOCOCCAL ARTHRITIS, LEFT WRIST
C4269532|T037|S02.651B|ICD10CM|FRACTURE OF ANGLE OF RIGHT MANDIBLE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF ANGLE OF RIGHT MANDIBLE, 7THB
C2895331|T037|M48.55XA|ICD10CM|COLLAPSED VERTEBRA, NOT ELSEWHERE CLASSIFIED, THORACOLUMBAR REGION, INITIAL ENCOUNTER FOR FRACTURE|COLLAPSED VERTEBRA, NEC, THORACOLUMBAR REGION, INIT
C2882828|T047|I70.435|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF OTHER PART OF FOOT|ATHSCL AUTOL VEIN BYPASS OF RIGHT LEG W ULCER OTH PRT FOOT
C2882826|T047|I70.434|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF HEEL AND MIDFOOT|ATHSCL AUTOL VEIN BYPASS OF R LEG W ULCER OF HEEL AND MIDFT
C2882824|T047|I70.433|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF ANKLE|ATHSCL AUTOL VEIN BYPASS OF THE RIGHT LEG W ULCER OF ANKLE
C2882823|T047|I70.432|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF CALF|ATHSCL AUTOL VEIN BYPASS OF THE RIGHT LEG W ULCER OF CALF
C2882822|T047|I70.431|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF THIGH|ATHSCL AUTOL VEIN BYPASS OF THE RIGHT LEG W ULCER OF THIGH
C2882830|T047|I70.439|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF UNSPECIFIED SITE|ATHSCL AUTOL VEIN BYPASS OF RIGHT LEG W ULCER OF UNSP SITE
C2882829|T047|I70.438|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF OTHER PART OF LOWER LEG|ATHSCL AUTOL VEIN BYPASS OF R LEG W ULCER OTH PRT LOW LEG
C2905788|T037|X81.8XXS|ICD10CM|INTENTIONAL SELF-HARM BY JUMPING OR LYING IN FRONT OF OTHER MOVING OBJECT, SEQUELA|SLF-HRM BY JUMP OR LYING IN FRONT OF MOVING OBJECT, SEQUELA
C0342571|T047|E34.4|DMDICD10|CONSTITUTIONAL TALL STATURE|KONSTITUTIONELLER HOCHWUCHS
C2874706|T048|F16.29|ICD10CM|HALLUCINOGEN DEPENDENCE WITH UNSPECIFIED HALLUCINOGEN-INDUCED DISORDER|HALLUCINOGEN DEPENDENCE W UNSP HALLUCINOGEN-INDUCED DISORDER
C0024586|T047|E34.0|DMDICD10|CARCINOID SYNDROME|KARZINOID-SYNDROM
C4237360|T048|F16.20|ICD10CM|HALLUCINOGEN DEPENDENCE, UNCOMPLICATED|PHENCYCLIDINE USE DISORDER, SEVERE
C4509075|T048|F16.21|ICD10CM|HALLUCINOGEN DEPENDENCE, IN REMISSION|OTHER HALLUCINOGEN USE DISORDER, SEVERE, IN SUSTAINED REMISSION
C2835312|T037|S22.042A|ICD10CM|UNSTABLE BURST FRACTURE OF FOURTH THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSTABLE BURST FRACTURE OF FOURTH THORACIC VERTEBRA, INIT
C4268272|T048|F16.24|ICD10CM|HALLUCINOGEN DEPENDENCE WITH HALLUCINOGEN-INDUCED MOOD DISORDER|PHENCYCLIDINE USE DISORDER, SEVERE, WITH PHENCYCLIDINE-INDUCED DEPRESSIVE DISORDER
C2857051|T037|S72.091A|ICD10CM|OTHER FRACTURE OF HEAD AND NECK OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF HEAD AND NECK OF RIGHT FEMUR, INIT
C2857053|T037|S72.091C|ICD10CM|OTHER FRACTURE OF HEAD AND NECK OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|OTH FX HEAD/NECK OF RIGHT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2857052|T037|S72.091B|ICD10CM|OTHER FRACTURE OF HEAD AND NECK OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|OTH FX HEAD/NECK OF RIGHT FEMUR, INIT FOR OPN FX TYPE I/2
C2889192|T047|M05.271|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF RIGHT ANK/FT
C2869756|T037|S98.011D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT FOOT AT ANKLE LEVEL, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMP OF RIGHT FOOT AT ANKLE LEVEL, SUBS
C2876192|T037|T32.41|ICD10CM|CORROSIONS INVOLVING 40-49% OF BODY SURFACE WITH 10-19% THIRD DEGREE CORROSION|CORROS 40-49% OF BODY SURFACE W 10-19% THIRD DEGREE CORROS
C2848393|T037|S58.012A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT ELBOW LEVEL, LEFT ARM, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION AT ELBOW LEVEL, LEFT ARM, INIT
C2885558|T037|T63.322A|ICD10CM|TOXIC EFFECT OF VENOM OF TARANTULA, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF TARANTULA, SELF-HARM, INIT
C2848395|T037|S58.012S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT ELBOW LEVEL, LEFT ARM, SEQUELA|COMPLETE TRAUMATIC AMP AT ELBOW LEVEL, LEFT ARM, SEQUELA
C2885560|T037|T63.322S|ICD10CM|TOXIC EFFECT OF VENOM OF TARANTULA, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF TARANTULA, SELF-HARM, SEQUELA
C2833264|T037|S12.130A|ICD10CM|UNSPECIFIED TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP TRAUM DISPL SPONDYLOLYSIS OF SECOND CERVCAL VERT, INIT
C2874691|T048|F16.183|ICD10CM|HALLUCINOGEN ABUSE WITH HALLUCINOGEN PERSISTING PERCEPTION DISORDER (FLASHBACKS)|HALLUCIGN ABUSE W HALLUCIGN PERSISTING PERCEPTION DISORDER
C2837647|T037|S32.058B|ICD10CM|OTHER FRACTURE OF FIFTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF FIFTH LUMBAR VERTEBRA, INIT FOR OPN FX
C2837646|T037|S32.058A|ICD10CM|OTHER FRACTURE OF FIFTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF FIFTH LUMBAR VERTEBRA, INIT FOR CLOS FX
C2901916|T047|M86.621|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, RIGHT  HUMERUS|OTHER CHRONIC OSTEOMYELITIS, RIGHT HUMERUS
C2874236|T047|E71.118|ICD10CM|OTHER BRANCHED-CHAIN ORGANIC ACIDURIAS|OTHER BRANCHED-CHAIN ORGANIC ACIDURIAS
C1260392|T047|E71.448|ICD10CM|OTHER SECONDARY CARNITINE DEFICIENCY|OTHER SECONDARY CARNITINE DEFICIENCY
C2834022|T037|S14.148D|ICD10CM|BROWN-SEQUARD SYNDROME AT C8 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|BROWN-SEQUARD SYNDROME AT C8, SUBS
C2833875|T037|S14.108D|ICD10CM|UNSPECIFIED INJURY AT C8 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY AT C8 LEVEL OF CERVICAL SPINAL CORD, SUBS ENCNTR
C3696376|T047||ICD10CM|3-METHYLGLUTACONIC ACIDURIA
C0268575|T047||ICD10CM|ISOVALERIC ACIDEMIA
C0265326|T047||ICD10CM|RUVALCABA-MYHRE-SMITH SYNDROME
C2858390|T037|S72.414B|ICD10CM|NONDISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP UNSP CONDYLE FX LOW END R FEMR, 7THB
C2858391|T037|S72.414C|ICD10CM|NONDISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP UNSP CONDYLE FX LOW END R FEMR, 7THC
C2858389|T037|S72.414A|ICD10CM|NONDISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP UNSP CONDYLE FX LOWER END OF RIGHT FEMUR, INIT
C2838085|T037|S32.426A|ICD10CM|NONDISPLACED FRACTURE OF POSTERIOR WALL OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF POSTERIOR WALL OF UNSP ACETABULUM, INIT
C2834023|T037|S14.148S|ICD10CM|BROWN-SEQUARD SYNDROME AT C8 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|BROWN-SEQUARD SYNDROME AT C8, SEQUELA
C4268098|T047|E11.3522|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, LEFT EYE|TYPE 2 DIAB W PROLIF DIAB RTNOP W TRCTN DTCH MACULA, L EYE
C4268099|T047|E11.3523|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, BILATERAL|TYPE 2 DIAB W PROLIF DIAB RTNOP WITH TRCTN DTCH MACULA, BI
C4268097|T047|E11.3521|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, RIGHT EYE|TYPE 2 DIAB W PROLIF DIAB RTNOP W TRCTN DTCH MACULA, R EYE
C2874246|T047|E71.4|ICD10CM|DISORDER OF CARNITINE METABOLISM, UNSPECIFIED|DISORDERS OF CARNITINE METABOLISM
C0342788|T047|E71.41|ICD10CM|PRIMARY CARNITINE DEFICIENCY|PRIMARY CARNITINE DEFICIENCY
C3875374|T047||ICD10CM|CARNITINE DEFICIENCY DUE TO INBORN ERRORS OF METABOLISM
C1260391|T046|E71.43|ICD10CM|IATROGENIC CARNITINE DEFICIENCY|IATROGENIC CARNITINE DEFICIENCY
C4268100|T047|E11.3529|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, UNSPECIFIED EYE|TYPE 2 DIAB W PROLIF DIAB RTNOP WITH TRCTN DTCH MACULA, UNSP
C0041806|T047|D89.9|DMDICD10|DISORDER INVOLVING THE IMMUNE MECHANISM, UNSPECIFIED|STOERUNG MIT BETEILIGUNG DES IMMUNSYSTEMS, NICHT NAEHER BEZEICHNET
C2976853|T047||ICD10CM|IMMUNE RECONSTITUTION SYNDROME
C2873857|T047|D89.1|ICD10CM|CRYOGLOBULINEMIA|IDIOPATHIC CRYOGLOBULINEMIA
C2833265|T037|S12.130B|ICD10CM|UNSPECIFIED TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP TRAUM DISPL SPONDYLOLYSIS OF 2ND CERVCAL VERT, 7THB
C0428981|T046|I49.2|DMDICD10|JUNCTIONAL PREMATURE DEPOLARIZATION|AV-JUNKTIONALE EXTRASYSTOLIE
C0221047|T047||ICD10CM|SICK SINUS SYNDROME
C2890747|T037|T84.310A|ICD10CM|BREAKDOWN (MECHANICAL) OF ELECTRONIC BONE STIMULATOR, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF ELECTRONIC BONE STIMULATOR, INIT
C2835211|T037|S22.018A|ICD10CM|OTHER FRACTURE OF FIRST THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF FIRST THORACIC VERTEBRA, INIT FOR CLOS FX
C4065471|T048|F34.81|ICD10CM|DISRUPTIVE MOOD DYSREGULATION DISORDER|DISRUPTIVE MOOD DYSREGULATION DISORDER
C4268303|T048|F34.89|ICD10CM|OTHER SPECIFIED PERSISTENT MOOD DISORDERS|OTHER SPECIFIED PERSISTENT MOOD DISORDERS
C0574027|T047||ICD10CM|ANEURYSM OF VERTEBRAL ARTERY
C0155744|T190|I72.4|DMDICD10|ANEURYSM OF ARTERY OF LOWER EXTREMITY|ANEURYSMA EINER ARTERIE DER UNTEREN EXTREMITAET
C4268547|T047|I72.5|ICD10CM|ANEURYSM OF OTHER PRECEREBRAL ARTERIES|ANEURYSM OF BASILAR ARTERY (TRUNK)
C0155742|T190|I72.2|DMDICD10|ANEURYSM OF RENAL ARTERY|ANEURYSMA DER NIERENARTERIE
C0162870|T190|I72.3|DMDICD10|ANEURYSM OF ILIAC ARTERY|ANEURYSMA DER A. ILIACA
C0865708|T190||ICD10CM|ANEURYSM OF CAROTID ARTERY
C0155741|T190|I72.1|DMDICD10|ANEURYSM OF ARTERY OF UPPER EXTREMITY|ANEURYSMA EINER ARTERIE DER OBEREN EXTREMITAET
C2896691|T046|M80.822A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, LEFT HUMERUS, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, L HUMERUS, INIT
C0002945|T190|I72.8|DMDICD10|ANEURYSM OF OTHER SPECIFIED ARTERIES|ANEURYSMA SONSTIGER NAEHER BEZEICHNETER ARTERIEN
C0002940|T190|I72.9|DMDICD10|ANEURYSM OF UNSPECIFIED SITE|ANEURYSMA NICHT NAEHER BEZEICHNETER LOKALISATION
C2835777|T037|S24.111D|ICD10CM|COMPLETE LESION AT T1 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION AT T1 LEVEL OF THORACIC SPINAL CORD, SUBS
C2835776|T037|S24.111A|ICD10CM|COMPLETE LESION AT T1 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION AT T1 LEVEL OF THORACIC SPINAL CORD, INIT
C2858679|T037|S72.443B|ICD10CM|DISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF LOW EPIPHY (SEPARATION) OF UNSP FEMR, 7THB
C2884286|T037|T53.5X2A|ICD10CM|TOXIC EFFECT OF CHLOROFLUOROCARBONS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CHLOROFLUOROCARBONS, SELF-HARM, INIT
C2858680|T037|S72.443C|ICD10CM|DISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF LOW EPIPHY (SEPARATION) OF UNSP FEMR, 7THC
C2885507|T037|T63.2X2A|ICD10CM|TOXIC EFFECT OF VENOM OF SCORPION, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF SCORPION, SELF-HARM, INIT
C2835778|T037|S24.111S|ICD10CM|COMPLETE LESION AT T1 LEVEL OF THORACIC SPINAL CORD, SEQUELA|COMPLETE LESION AT T1 LEVEL OF THORACIC SPINAL CORD, SEQUELA
C2884288|T037|T53.5X2S|ICD10CM|TOXIC EFFECT OF CHLOROFLUOROCARBONS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CHLOROFLUOROCARBONS, SELF-HARM, SEQUELA
C2900975|T046|M84.445A|ICD10CM|PATHOLOGICAL FRACTURE, LEFT FINGER(S), INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, LEFT FINGER(S), INIT FOR FX
C2900918|T046|M84.432A|ICD10CM|PATHOLOGICAL FRACTURE, LEFT ULNA, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, LEFT ULNA, INIT ENCNTR FOR FRACTURE
C2902086|T046|M87.32|ICD10CM|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED HUMERUS|OTHER SECONDARY OSTEONECROSIS, HUMERUS
C2910918|T033|Z48.24|ICD10CM|ENCOUNTER FOR AFTERCARE FOLLOWING LUNG TRANSPLANT|ENCOUNTER FOR AFTERCARE FOLLOWING LUNG TRANSPLANT
C2902084|T046|M87.321|ICD10CM|OTHER SECONDARY OSTEONECROSIS, RIGHT HUMERUS|OTHER SECONDARY OSTEONECROSIS, RIGHT HUMERUS
C2902085|T046|M87.322|ICD10CM|OTHER SECONDARY OSTEONECROSIS, LEFT HUMERUS|OTHER SECONDARY OSTEONECROSIS, LEFT HUMERUS
C2882719|T047|I70.239|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF RIGHT LEG WITH ULCERATION OF UNSPECIFIED SITE|ATHSCL NATIVE ARTERIES OF RIGHT LEG W ULCER OF UNSP SITE
C2882718|T047|I70.238|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF RIGHT LEG WITH ULCERATION OF OTHER PART OF LOWER RIGHT LEG|ATHSCL NATV ART OF RIGHT LEG W ULCER OTH PRT LOWER RIGHT LEG
C2882717|T047|I70.235|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF RIGHT LEG WITH ULCERATION OF OTHER PART OF FOOT|ATHSCL NATIVE ARTERIES OF RIGHT LEG W ULCER OTH PRT FOOT
C2882715|T047|I70.234|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF RIGHT LEG WITH ULCERATION OF HEEL AND MIDFOOT|ATHSCL NATIVE ART OF RIGHT LEG W ULCER OF HEEL AND MIDFOOT
C2882711|T047|I70.231|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF RIGHT LEG WITH ULCERATION OF THIGH|ATHSCL NATIVE ARTERIES OF RIGHT LEG W ULCERATION OF THIGH
C2882713|T047|I70.233|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF RIGHT LEG WITH ULCERATION OF ANKLE|ATHSCL NATIVE ARTERIES OF RIGHT LEG W ULCERATION OF ANKLE
C2882712|T047|I70.232|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF RIGHT LEG WITH ULCERATION OF CALF|ATHSCL NATIVE ARTERIES OF RIGHT LEG W ULCERATION OF CALF
C2874064|T047|E10.628|ICD10CM|TYPE 1 DIABETES MELLITUS WITH OTHER SKIN COMPLICATIONS|TYPE 1 DIABETES MELLITUS WITH OTHER SKIN COMPLICATIONS
C2887771|T047|K50.80|ICD10CM|CROHN'S DISEASE OF BOTH SMALL AND LARGE INTESTINE WITHOUT COMPLICATIONS|CROHN'S DISEASE OF BOTH SMALL AND LG INT W/O COMPLICATIONS
C2910917|T033|Z48.23|ICD10CM|ENCOUNTER FOR AFTERCARE FOLLOWING LIVER TRANSPLANT|ENCOUNTER FOR AFTERCARE FOLLOWING LIVER TRANSPLANT
C2890015|T037|T82.514A|ICD10CM|BREAKDOWN (MECHANICAL) OF INFUSION CATHETER, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF INFUSION CATHETER, INIT ENCNTR
C2874061|T047|E10.620|ICD10CM|TYPE 1 DIABETES MELLITUS WITH DIABETIC DERMATITIS|TYPE 1 DIABETES MELLITUS WITH DIABETIC DERMATITIS
C2874062|T047|E10.621|ICD10CM|TYPE 1 DIABETES MELLITUS WITH FOOT ULCER|TYPE 1 DIABETES MELLITUS WITH FOOT ULCER
C2874063|T047|E10.622|ICD10CM|TYPE 1 DIABETES MELLITUS WITH OTHER SKIN ULCER|TYPE 1 DIABETES MELLITUS WITH OTHER SKIN ULCER
C2858904|T037|S72.464C|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP SUPRCNDL FX W INTRCNDL EXTN LOW END R FEMR, 7THC
C2858560|T037|S72.432B|ICD10CM|DISPLACED FRACTURE OF MEDIAL CONDYLE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF MED CONDYLE OF L FEMUR, INIT FOR OPN FX TYPE I/2
C2858561|T037|S72.432C|ICD10CM|DISPLACED FRACTURE OF MEDIAL CONDYLE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF MED CONDYLE OF L FEMR, 7THC
C2834064|T037|S14.159A|ICD10CM|OTHER INCOMPLETE LESION AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|OTH INCMPL LESION AT UNSP LEVEL OF CERV SPINAL CORD, INIT
C2860010|T037|S78.121A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN RIGHT HIP AND KNEE, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP AT LEVEL BETW RIGHT HIP AND KNEE, INIT
C2860011|T037|S78.121D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN RIGHT HIP AND KNEE, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMP AT LEVEL BETW RIGHT HIP AND KNEE, SUBS
C4267974|T047|E09.3491|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|DRUG/CHEM DIAB WITH SEVERE NONP RTNOP W/O MCLR EDEMA, R EYE
C4267976|T047|E09.3493|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|DRUG/CHEM DIAB WITH SEVERE NONP RTNOP WITHOUT MCLR EDEMA, BI
C4267975|T047|E09.3492|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|DRUG/CHEM DIAB WITH SEVERE NONP RTNOP W/O MCLR EDEMA, L EYE
C4267977|T047|E09.3499|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|DRUG/CHEM DIAB WITH SEVERE NONP RTNOP W/O MCLR EDEMA, UNSP
C2889950|T037|T82.339A|ICD10CM|LEAKAGE OF UNSPECIFIED VASCULAR GRAFT, INITIAL ENCOUNTER|LEAKAGE OF UNSPECIFIED VASCULAR GRAFT, INITIAL ENCOUNTER
C2856011|T037|S68.612S|ICD10CM|COMPLETE TRAUMATIC TRANSPHALANGEAL AMPUTATION OF RIGHT MIDDLE FINGER, SEQUELA|COMPLETE TRAUMATIC TRNSPHAL AMP OF R MID FINGER, SEQUELA
C2832066|T037|S06.303A|ICD10CM|UNSPECIFIED FOCAL TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|UNSP FOCAL TBI W LOC OF 1-5 HRS 59 MIN, INIT
C2888394|T047||ICD10CM|PRESSURE ULCER OF LEFT HIP, UNSTAGEABLE
C2901191|T046|M84.532A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, LEFT ULNA, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, LEFT ULNA, INIT
C2901234|T046|M84.549A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, UNSPECIFIED HAND, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, UNSP HAND, INIT
C2832068|T037|S06.303S|ICD10CM|UNSPECIFIED FOCAL TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, SEQUELA|UNSP FOCAL TBI W LOC OF 1-5 HRS 59 MIN, SEQUELA
C2877715|T037|T40.602S|ICD10CM|POISONING BY UNSPECIFIED NARCOTICS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY UNSP NARCOTICS, INTENTIONAL SELF-HARM, SEQUELA
C2896485|T046|M80.011A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, RIGHT SHOULDER, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, R SHOULDER, INIT
C2884819|T037|T58.92XS|ICD10CM|TOXIC EFFECT OF CARBON MONOXIDE FROM UNSPECIFIED SOURCE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CARB MONX FROM UNSP SOURCE, SLF-HRM, SEQUELA
C2890805|T037|T84.51XA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL RIGHT HIP PROSTHESIS, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INTERNAL RIGHT HIP PROSTH, INIT
C2887313|T047|I87.339|ICD10CM|CHRONIC VENOUS HYPERTENSION (IDIOPATHIC) WITH ULCER AND INFLAMMATION OF UNSPECIFIED LOWER EXTREMITY|CHRONIC VENOUS HTN W ULCER AND INFLAM OF UNSP LOW EXTRM
C2888681|T047|L97.309|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED ANKLE WITH UNSPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF UNSP ANKLE WITH UNSP SEVERITY
C2884817|T037|T58.92XA|ICD10CM|TOXIC EFFECT OF CARBON MONOXIDE FROM UNSPECIFIED SOURCE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CARB MONX FROM UNSP SOURCE, SELF-HARM, INIT
C4509295|T047|L97.308|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED ANKLE WITH OTHER SPECIFIED SEVERITY|NON-PRS CHRONIC ULCER OF UNSPECIFIED ANKLE WITH OTH SEVERITY
C2877279|T037|T38.902A|ICD10CM|POISONING BY UNSPECIFIED HORMONE ANTAGONISTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY UNSP HORMONE ANTAGONISTS, SELF-HARM, INIT
C2889058|T047|M02.331|ICD10CM|REITER'S DISEASE, RIGHT WRIST|REITER'S DISEASE, RIGHT WRIST
C2901971|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF RIGHT FIBULA
C0494293|T047|E13.9|DMDICD10|OTHER SPECIFIED DIABETES MELLITUS WITHOUT COMPLICATIONS|SONSTIGER NAEHER BEZEICHNETER DIABETES MELLITUS: OHNE KOMPLIKATIONEN
C2889059|T047|M02.332|ICD10CM|REITER'S DISEASE, LEFT WRIST|REITER'S DISEASE, LEFT WRIST
C2874224|T047|E64.0|ICD10CM|SEQUELAE OF PROTEIN-CALORIE MALNUTRITION|SEQUELAE OF PROTEIN-CALORIE MALNUTRITION
C2889060|T047|M02.339|ICD10CM|REITER'S DISEASE, UNSPECIFIED WRIST|REITER'S DISEASE, UNSPECIFIED WRIST
C2888375|T047|L89.209|ICD10CM|PRESSURE ULCER OF UNSPECIFIED HIP, UNSPECIFIED STAGE|PRESSURE ULCER OF UNSPECIFIED HIP, UNSPECIFIED STAGE
C2877948|T037|T41.292S|ICD10CM|POISONING BY OTHER GENERAL ANESTHETICS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH GENERAL ANESTHETICS, SELF-HARM, SEQUELA
C2888369|T047|L89.203|ICD10CM|PRESSURE ULCER OF UNSPECIFIED HIP, STAGE 3|PRESSURE ULCER OF UNSPECIFIED HIP, STAGE 3
C2888366|T047|L89.202|ICD10CM|PRESSURE ULCER OF UNSPECIFIED HIP, STAGE 2|PRESSURE ULCER OF UNSPECIFIED HIP, STAGE 2
C2888363|T047|L89.201|ICD10CM|PRESSURE ULCER OF UNSPECIFIED HIP, STAGE 1|PRESSURE ULCER OF UNSPECIFIED HIP, STAGE 1
C2888360|T047|L89.200|ICD10CM|PRESSURE ULCER OF UNSPECIFIED HIP, UNSTAGEABLE|PRESSURE ULCER OF UNSPECIFIED HIP, UNSTAGEABLE
C2888372|T047|L89.204|ICD10CM|PRESSURE ULCER OF UNSPECIFIED HIP, STAGE 4|PRESSURE ULCER OF UNSPECIFIED HIP, STAGE 4
C2882462|T047|I69.049|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING UNSPECIFIED SIDE|MONOPLG LOW LMB FOLLOWING NTRM SUBARACH HEMOR AFF UNSP SIDE
C2882458|T047|I69.041|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING RIGHT DOMINANT SIDE|MONOPLG LOW LMB FOL NTRM SUBARACH HEMOR AFF RIGHT DOM SIDE
C2882459|T047|I69.042|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING LEFT DOMINANT SIDE|MONOPLG LOW LMB FOL NTRM SUBARACH HEMOR AFF LEFT DOM SIDE
C2882460|T047|I69.043|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING RIGHT NON-DOMINANT SIDE|MONOPLG LOW LMB FOL NTRM SUBARACH HEMOR AFF R NONDOM SIDE
C2882461|T047|I69.044|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING LEFT NON-DOMINANT SIDE|MONOPLG LOW LMB FOL NTRM SUBARACH HEMOR AFF LEFT NONDOM SIDE
C2838300|T037|S32.476A|ICD10CM|NONDISPLACED FRACTURE OF MEDIAL WALL OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF MEDIAL WALL OF UNSP ACETABULUM, INIT
C2888679|T047|L97.303|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED ANKLE WITH NECROSIS OF MUSCLE|NON-PRS CHRONIC ULCER OF UNSP ANKLE W NECROSIS OF MUSCLE
C2876547|T037|T36.0X2S|ICD10CM|POISONING BY PENICILLINS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY PENICILLINS, INTENTIONAL SELF-HARM, SEQUELA
C2711480|T047||ICD10CM|CHRONIC DIASTOLIC (CONGESTIVE) HEART FAILURE
C2732749|T047||ICD10CM|ACUTE ON CHRONIC DIASTOLIC (CONGESTIVE) HEART FAILURE
C1135196|T047|I50.30|ICD10CM|UNSPECIFIED DIASTOLIC (CONGESTIVE) HEART FAILURE|UNSPECIFIED DIASTOLIC (CONGESTIVE) HEART FAILURE
C2215111|T047||ICD10CM|ACUTE DIASTOLIC (CONGESTIVE) HEART FAILURE
C2889994|T037|T82.49XA|ICD10CM|OTHER COMPLICATION OF VASCULAR DIALYSIS CATHETER, INITIAL ENCOUNTER|OTH COMPLICATION OF VASCULAR DIALYSIS CATHETER, INIT ENCNTR
C2905750|T037|X78.0XXA|ICD10CM|INTENTIONAL SELF-HARM BY SHARP GLASS, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY SHARP GLASS, INITIAL ENCOUNTER
C2884352|T037|T54.0X2S|ICD10CM|TOXIC EFFECT OF PHENOL AND PHENOL HOMOLOGUES, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF PHENOL AND PHENOL HOMOLOG, SLF-HRM, SEQUELA
C2875095|T047|G40.211|ICD10CM|LOCALIZATION-RELATED (FOCAL) (PARTIAL) SYMPTOMATIC EPILEPSY AND EPILEPTIC SYNDROMES WITH COMPLEX PARTIAL SEIZURES, INTRACTABLE, WITH STATUS EPILEPTICUS|LOCAL-REL SYMPTC EPI W CMPLX PARTIAL SEIZ, NTRCT, W STAT EPI
C2367455|T191||ICD10CM|ACUTE MEGAKARYOBLASTIC LEUKEMIA, IN RELAPSE
C0153914|T191||ICD10AM|ACUTE MEGAKARYOBLASTIC LEUKEMIA, IN REMISSION
C2861634|T191|C94.20|ICD10CM|ACUTE MEGAKARYOBLASTIC LEUKEMIA NOT HAVING ACHIEVED REMISSION|ACUTE MEGAKARYOBLASTIC LEUKEMIA WITH FAILED REMISSION
C2889996|T037|T82.49XS|ICD10CM|OTHER COMPLICATION OF VASCULAR DIALYSIS CATHETER, SEQUELA|OTHER COMPLICATION OF VASCULAR DIALYSIS CATHETER, SEQUELA
C2884350|T037|T54.0X2A|ICD10CM|TOXIC EFFECT OF PHENOL AND PHENOL HOMOLOGUES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF PHENOL AND PHENOL HOMOLOG, SELF-HARM, INIT
C2853917|T191|C83.38|ICD10CM|DIFFUSE LARGE B-CELL LYMPHOMA, LYMPH NODES OF MULTIPLE SITES|DIFFUSE LARGE B-CELL LYMPHOMA, LYMPH NODES OF MULTIPLE SITES
C3647864|T191|C83.39|ICD10CM|DIFFUSE LARGE B-CELL LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES|DIFFUSE LARGE B-CELL LYMPHOMA, EXTRNOD AND SOLID ORGAN SITES
C2893630|T047|M12.012|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], LEFT SHOULDER|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], LEFT SHOULDER
C2853914|T191|C83.34|ICD10CM|DIFFUSE LARGE B-CELL LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB|DIFFUSE LARGE B-CELL LYMPH, NODES OF AXILLA AND UPPER LIMB
C2853915|T191|C83.35|ICD10CM|DIFFUSE LARGE B-CELL LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|DIFFUS LARGE B-CELL LYMPH, NODES OF ING RGN AND LOWER LIMB
C2853916|T191|C83.36|ICD10CM|DIFFUSE LARGE B-CELL LYMPHOMA, INTRAPELVIC LYMPH NODES|DIFFUSE LARGE B-CELL LYMPHOMA, INTRAPELVIC LYMPH NODES
C2018774|T191||ICD10CM|DIFFUSE LARGE B-CELL LYMPHOMA, SPLEEN
C2853910|T191|C83.30|ICD10CM|DIFFUSE LARGE B-CELL LYMPHOMA, UNSPECIFIED SITE|DIFFUSE LARGE B-CELL LYMPHOMA, UNSPECIFIED SITE
C2853911|T191|C83.31|ICD10CM|DIFFUSE LARGE B-CELL LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK|DIFFUSE LARGE B-CELL LYMPHOMA, NODES OF HEAD, FACE, AND NECK
C2853912|T191|C83.32|ICD10CM|DIFFUSE LARGE B-CELL LYMPHOMA, INTRATHORACIC LYMPH NODES|DIFFUSE LARGE B-CELL LYMPHOMA, INTRATHORACIC LYMPH NODES
C2853913|T191|C83.33|ICD10CM|DIFFUSE LARGE B-CELL LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES|DIFFUSE LARGE B-CELL LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES
C2875096|T047|G40.219|ICD10CM|LOCALIZATION-RELATED (FOCAL) (PARTIAL) SYMPTOMATIC EPILEPSY AND EPILEPTIC SYNDROMES WITH COMPLEX PARTIAL SEIZURES, INTRACTABLE, WITHOUT STATUS EPILEPTICUS|LOCAL-REL SYMPTC EPI W CMPLX PART SEIZ, NTRCT, W/O STAT EPI
C4270459|T046|T85.111A|ICD10CM|BREAKDOWN (MECHANICAL) OF IMPLANTED ELECTRONIC NEUROSTIMULATOR OF PERIPHERAL NERVE ELECTRODE (LEAD), INITIAL ENCOUNTER|BREAKDOWN OF IMPLNT ELEC NSTIM OF PRPH NRV LEAD, INIT
C2905751|T037|X78.0XXD|ICD10CM|INTENTIONAL SELF-HARM BY SHARP GLASS, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY SHARP GLASS, SUBSEQUENT ENCOUNTER
C2875162|T047|G43.509|ICD10CM|PERSISTENT MIGRAINE AURA WITHOUT CEREBRAL INFARCTION, NOT INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|PERST MIGRN AURA W/O CEREB INFRC, NOT NTRCT, W/O STAT MIGR
C2875161|T047|G43.501|ICD10CM|PERSISTENT MIGRAINE AURA WITHOUT CEREBRAL INFARCTION, NOT INTRACTABLE, WITH STATUS MIGRAINOSUS|PERST MIGRAINE AURA W/O CEREB INFRC, NOT NTRCT, W STAT MIGR
C2882185|T047|I25.721|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS ARTERY CORONARY ARTERY BYPASS GRAFT(S) WITH ANGINA PECTORIS WITH DOCUMENTED SPASM|ATHSCL AUTOLOGOUS ARTERY CABG W ANG PCTRS W DOCUMENTED SPASM
C4270569|T046|T85.730A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO VENTRICULAR INTRACRANIAL (COMMUNICATING) SHUNT, INITIAL ENCOUNTER|I/I REACT D/T VENTRICULAR INTRACRANIAL SHUNT, INIT
C2843279|T037|S48.019S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT UNSPECIFIED SHOULDER JOINT, SEQUELA|COMPLETE TRAUMATIC AMPUTATION AT UNSP SHOULDER JT, SEQUELA
C2837826|T037|S32.311B|ICD10CM|DISPLACED AVULSION FRACTURE OF RIGHT ILIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISPLACED AVULSION FRACTURE OF RIGHT ILIUM, INIT FOR OPN FX
C2890397|T037|T83.9XXA|ICD10CM|UNSPECIFIED COMPLICATION OF GENITOURINARY PROSTHETIC DEVICE, IMPLANT AND GRAFT, INITIAL ENCOUNTER|UNSP COMPLICATION OF GENITOURINARY PROSTH DEV/GRFT, INIT
C2889613|T047|M08.849|ICD10CM|OTHER JUVENILE ARTHRITIS, UNSPECIFIED HAND|OTHER JUVENILE ARTHRITIS, UNSPECIFIED HAND
C4509340|T047|L98.418|ICD10CM|NON-PRESSURE CHRONIC ULCER OF BUTTOCK WITH OTHER SPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF BUTTOCK WITH OTH SEVERITY
C2888778|T047|L98.419|ICD10CM|NON-PRESSURE CHRONIC ULCER OF BUTTOCK WITH UNSPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF BUTTOCK WITH UNSP SEVERITY
C2882910|T047|I70.592|ICD10CM|OTHER ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, LEFT LEG|OTH ATHSCL NONAUT BIO BYPASS OF THE EXTREMITIES, LEFT LEG
C2882911|T047|I70.593|ICD10CM|OTHER ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, BILATERAL LEGS|OTH ATHSCL NONAUT BIO BYPASS OF THE EXTRM, BILATERAL LEGS
C2883075|T047|I80.239|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF UNSPECIFIED TIBIAL VEIN|PHLEBITIS AND THROMBOPHLEBITIS OF UNSPECIFIED TIBIAL VEIN
C2882912|T047|I70.598|ICD10CM|OTHER ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, OTHER EXTREMITY|OTH ATHSCL NONAUT BIO BYPASS OF THE EXTRM, OTH EXTREMITY
C2888774|T047|L98.411|ICD10CM|NON-PRESSURE CHRONIC ULCER OF BUTTOCK LIMITED TO BREAKDOWN OF SKIN|NON-PRESSURE CHRONIC ULCER OF BUTTOCK LIMITED TO BRKDWN SKIN
C2888775|T047||ICD10CM|NON-PRESSURE CHRONIC ULCER OF BUTTOCK WITH FAT LAYER EXPOSED
C2888776|T047|L98.413|ICD10CM|NON-PRESSURE CHRONIC ULCER OF BUTTOCK WITH NECROSIS OF MUSCLE|NON-PRESSURE CHRONIC ULCER OF BUTTOCK W NECROSIS OF MUSCLE
C2888777|T047||ICD10CM|NON-PRESSURE CHRONIC ULCER OF BUTTOCK WITH NECROSIS OF BONE
C4509338|T047|L98.415|ICD10CM|NON-PRESSURE CHRONIC ULCER OF BUTTOCK WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULCER OF BUTTOCK WITH MSL INVL W/O EVD OF NECR
C4509339|T047|L98.416|ICD10CM|NON-PRESSURE CHRONIC ULCER OF BUTTOCK WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULCER OF BUTTOCK WITH BONE INVL W/O EVD OF NECR
C2883072|T047|I80.231|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF RIGHT TIBIAL VEIN|PHLEBITIS AND THROMBOPHLEBITIS OF RIGHT TIBIAL VEIN
C2889555|T047|M08.221|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, RIGHT ELBOW|JUVENILE RHEUMATOID ARTHRITIS W SYSTEMIC ONSET, RIGHT ELBOW
C2889556|T047|M08.222|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, LEFT ELBOW|JUVENILE RHEUMATOID ARTHRITIS W SYSTEMIC ONSET, LEFT ELBOW
C2878976|T037|T44.902S|ICD10CM|POISONING BY UNSPECIFIED DRUGS PRIMARILY AFFECTING THE AUTONOMIC NERVOUS SYSTEM, INTENTIONAL SELF-HARM, SEQUELA|POISN BY UNSP DRUGS AFF THE AUTONM NRV SYS, SLF-HRM, SEQUELA
C2889554|T047|M08.22|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, UNSPECIFIED ELBOW|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, ELBOW
C2857222|T037|S72.115A|ICD10CM|NONDISPLACED FRACTURE OF GREATER TROCHANTER OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF GREATER TROCHANTER OF LEFT FEMUR, INIT
C0221227|T047|J43.2|DMDICD10|CENTRILOBULAR EMPHYSEMA|ZENTRILOBULAERES EMPHYSEM
C0264393|T047|J43.1|DMDICD10|PANLOBULAR EMPHYSEMA|PANLOBULAERES EMPHYSEM
C2887442|T047|J43.0|ICD10CM|UNILATERAL PULMONARY EMPHYSEMA [MACLEOD'S SYNDROME]|UNILATERAL PULMONARY EMPHYSEMA [MACLEOD'S SYNDROME]
C2887444|T047|J43.9|ICD10CM|EMPHYSEMA, UNSPECIFIED|VESICULAR EMPHYSEMA (LUNG)(PULMONARY)
C0029607|T047|J43.8|DMDICD10|OTHER EMPHYSEMA|SONSTIGES EMPHYSEM
C0837456|T047||ICD10CM|OTHER REACTIVE ARTHROPATHIES, UNSPECIFIED SITE
C2837868|T037|S32.391A|ICD10CM|OTHER FRACTURE OF RIGHT ILIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF RIGHT ILIUM, INIT ENCNTR FOR CLOSED FRACTURE
C2889104|T047|M02.88|ICD10CM|OTHER REACTIVE ARTHROPATHIES, VERTEBRAE|OTHER REACTIVE ARTHROPATHIES, VERTEBRAE
C0837456|T047|M02.89|ICD10AM|OTHER REACTIVE ARTHROPATHIES, MULTIPLE SITES|OTHER REACTIVE ARTHROPATHIES, SITE UNSPECIFIED
C2833899|T037|S14.115D|ICD10CM|COMPLETE LESION AT C5 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION AT C5 LEVEL OF CERVICAL SPINAL CORD, SUBS
C2857325|T037|S72.125A|ICD10CM|NONDISPLACED FRACTURE OF LESSER TROCHANTER OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF LESSER TROCHANTER OF LEFT FEMUR, INIT
C2857327|T037|S72.125C|ICD10CM|NONDISPLACED FRACTURE OF LESSER TROCHANTER OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF LESS TROCHANTER OF L FEMR, 7THC
C2857326|T037|S72.125B|ICD10CM|NONDISPLACED FRACTURE OF LESSER TROCHANTER OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF LESS TROCHANTER OF L FEMR, 7THB
C2833970|T037|S14.134S|ICD10CM|ANTERIOR CORD SYNDROME AT C4 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|ANTERIOR CORD SYNDROME AT C4, SEQUELA
C0837021|T047|E11.00|ICD10CM|TYPE 2 DIABETES MELLITUS WITH HYPEROSMOLARITY WITHOUT NONKETOTIC HYPERGLYCEMIC-HYPEROSMOLAR COMA (NKHHC)|TYPE 2 DIAB W HYPROSM W/O NONKET HYPRGLY-HYPROS COMA (NKHHC)
C0837022|T047|E11.01|ICD10CM|TYPE 2 DIABETES MELLITUS WITH HYPEROSMOLARITY WITH COMA|TYPE 2 DIABETES MELLITUS WITH HYPEROSMOLARITY WITH COMA
C2883035|T047|I73.01|ICD10CM|RAYNAUD'S SYNDROME WITH GANGRENE|RAYNAUD'S SYNDROME WITH GANGRENE
C2833969|T037|S14.134D|ICD10CM|ANTERIOR CORD SYNDROME AT C4 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|ANTERIOR CORD SYNDROME AT C4, SUBS
C2833968|T037|S14.134A|ICD10CM|ANTERIOR CORD SYNDROME AT C4 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|ANTERIOR CORD SYNDROME AT C4, INIT
C2856741|T037|S72.034A|ICD10CM|NONDISPLACED MIDCERVICAL FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED MIDCERVICAL FRACTURE OF RIGHT FEMUR, INIT
C2856742|T037|S72.034B|ICD10CM|NONDISPLACED MIDCERVICAL FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP MIDCERVICAL FX RIGHT FEMUR, INIT FOR OPN FX TYPE I/2
C2856743|T037|S72.034C|ICD10CM|NONDISPLACED MIDCERVICAL FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP MIDCERVICAL FX R FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2869842|T037|S98.219A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF TWO OR MORE UNSPECIFIED LESSER TOES, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMP OF TWO OR MORE UNSP LESSER TOES, INIT
C2873778|T047|D61.01|ICD10CM|CONSTITUTIONAL (PURE) RED BLOOD CELL APLASIA|CONSTITUTIONAL (PURE) RED BLOOD CELL APLASIA
C0496933|T191|D42.0|DMDICD10|NEOPLASM OF UNCERTAIN BEHAVIOR OF CEREBRAL MENINGES|NEUBILDUNG UNSICHEREN ODER UNBEKANNTEN VERHALTENS: HIRNHAEUTE
C0496934|T191|D42.1|DMDICD10|NEOPLASM OF UNCERTAIN BEHAVIOR OF SPINAL MENINGES|NEUBILDUNG UNSICHEREN ODER UNBEKANNTEN VERHALTENS: RUECKENMARKHAEUTE
C3648009|T191||ICD10CM|CUTANEOUS FOLLICLE CENTER LYMPHOMA, INTRAPELVIC LYMPH NODES
C4269546|T037|S02.670B|ICD10CM|FRACTURE OF ALVEOLUS OF MANDIBLE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF ALVEOLUS OF MANDIBLE, UNSPECIFIED SIDE, 7THB
C4269545|T037|S02.670A|ICD10CM|FRACTURE OF ALVEOLUS OF MANDIBLE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF ALVEOLUS OF MANDIBLE, UNSPECIFIED SIDE, INIT
C2845985|T191|C7B.8|ICD10CM|OTHER SECONDARY NEUROENDOCRINE TUMORS|OTHER SECONDARY NEUROENDOCRINE TUMORS
C2877048|T037|T38.2X2S|ICD10CM|POISONING BY ANTITHYROID DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ANTITHYROID DRUGS, SELF-HARM, SEQUELA
C2856638|T037|S72.024B|ICD10CM|NONDISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF EPIPHY (SEPARATION) (UPPER) OF R FEMR, 7THB
C2712933|T191||ICD10CM|SECONDARY MERKEL CELL CARCINOMA
C0003869|T047|M00|DMDICD10|PYOGENIC ARTHRITIS, UNSPECIFIED|EITRIGE ARTHRITIS
C0839958|T047|M86.30|ICD10AM|CHRONIC MULTIFOCAL OSTEOMYELITIS, UNSPECIFIED SITE|CHRONIC MULTIFOCAL OSTEOMYELITIS, MULTIPLE SITES
C2902000|T046|M87.138|ICD10CM|OSTEONECROSIS DUE TO DRUGS OF LEFT CARPUS|OSTEONECROSIS DUE TO DRUGS OF LEFT CARPUS
C2902001|T046|M87.139|ICD10CM|OSTEONECROSIS DUE TO DRUGS OF UNSPECIFIED CARPUS|OSTEONECROSIS DUE TO DRUGS OF UNSPECIFIED CARPUS
C2901996|T046|M87.134|ICD10CM|OSTEONECROSIS DUE TO DRUGS OF RIGHT ULNA|OSTEONECROSIS DUE TO DRUGS OF RIGHT ULNA
C2901997|T046|M87.135|ICD10CM|OSTEONECROSIS DUE TO DRUGS OF LEFT ULNA|OSTEONECROSIS DUE TO DRUGS OF LEFT ULNA
C0839958|T047|M86.39|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, MULTIPLE SITES|CHRONIC MULTIFOCAL OSTEOMYELITIS, MULTIPLE SITES
C0839966|T047|M86.38|ICD10AM|CHRONIC MULTIFOCAL OSTEOMYELITIS, OTHER SITE|CHRONIC MULTIFOCAL OSTEOMYELITIS, OTHER SITE
C2901993|T046|M87.131|ICD10CM|OSTEONECROSIS DUE TO DRUGS OF RIGHT RADIUS|OSTEONECROSIS DUE TO DRUGS OF RIGHT RADIUS
C2901994|T046|M87.132|ICD10CM|OSTEONECROSIS DUE TO DRUGS OF LEFT RADIUS|OSTEONECROSIS DUE TO DRUGS OF LEFT RADIUS
C2901995|T046|M87.133|ICD10CM|OSTEONECROSIS DUE TO DRUGS OF UNSPECIFIED RADIUS|OSTEONECROSIS DUE TO DRUGS OF UNSPECIFIED RADIUS
C2889202|T047|M05.319|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP SHOULDER
C2879308|T037|T45.7X2A|ICD10CM|POISONING BY ANTICOAGULANT ANTAGONISTS, VITAMIN K AND OTHER COAGULANTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY ANTICOAG ANTAG, VIT K AND OTH COAG, SLF-HRM, INIT
C2889201|T047|M05.312|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT SHOULDER|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF L SHOULDER
C2889200|T047|M05.311|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT SHOULDER|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF R SHOULDER
C2883661|T037|T50.5X2S|ICD10CM|POISONING BY APPETITE DEPRESSANTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY APPETITE DEPRESSANTS, SELF-HARM, SEQUELA
C2848458|T037|S58.922A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT FOREARM, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF L FOREARM, LEVEL UNSP, INIT
C2887812|T047|K51.40|ICD10CM|INFLAMMATORY POLYPS OF COLON WITHOUT COMPLICATIONS|INFLAMMATORY POLYPS OF COLON WITHOUT COMPLICATIONS
C4270185|T046|T83.011A|ICD10CM|BREAKDOWN (MECHANICAL) OF INDWELLING URETHRAL CATHETER, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF INDWELLING URETHRAL CATHETER, INIT
C2889089|T047|M02.839|ICD10CM|OTHER REACTIVE ARTHROPATHIES, UNSPECIFIED WRIST|OTHER REACTIVE ARTHROPATHIES, UNSPECIFIED WRIST
C2889088|T047|M02.832|ICD10CM|OTHER REACTIVE ARTHROPATHIES, LEFT WRIST|OTHER REACTIVE ARTHROPATHIES, LEFT WRIST
C2889087|T047|M02.831|ICD10CM|OTHER REACTIVE ARTHROPATHIES, RIGHT WRIST|OTHER REACTIVE ARTHROPATHIES, RIGHT WRIST
C2858729|T037|S72.446A|ICD10CM|NONDISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF LOWER EPIPHY (SEPARATION) OF UNSP FEMUR, INIT
C2853894|T191|C83.10|ICD10CM|MANTLE CELL LYMPHOMA, UNSPECIFIED SITE|MANTLE CELL LYMPHOMA, UNSPECIFIED SITE
C2858731|T037|S72.446C|ICD10CM|NONDISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF LOW EPIPHY (SEPARATION) OF UNSP FEMR, 7THC
C2858730|T037|S72.446B|ICD10CM|NONDISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF LOW EPIPHY (SEPARATION) OF UNSP FEMR, 7THB
C2838641|T037|S34.111A|ICD10CM|COMPLETE LESION OF L1 LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION OF L1 LEVEL OF LUMBAR SPINAL CORD, INIT
C2838642|T037|S34.111D|ICD10CM|COMPLETE LESION OF L1 LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION OF L1 LEVEL OF LUMBAR SPINAL CORD, SUBS
C1386301|T047||ICD10CM|OTHER SPECIFIED METABOLIC DISORDERS
C2878660|T037|T43.692A|ICD10CM|POISONING BY OTHER PSYCHOSTIMULANTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH PSYCHOSTIMULANTS, SELF-HARM, INIT
C2861586|T191|C92.20|ICD10CM|ATYPICAL CHRONIC MYELOID LEUKEMIA, BCR/ABL-NEGATIVE, NOT HAVING ACHIEVED REMISSION|ATYP CHRONIC MYELOID LEUK, BCR/ABL-NEG, NOT ACHIEVE REMIS
C2845883|T191|C63.02|ICD10CM|MALIGNANT NEOPLASM OF LEFT EPIDIDYMIS|MALIGNANT NEOPLASM OF LEFT EPIDIDYMIS
C2845882|T191|C63.01|ICD10CM|MALIGNANT NEOPLASM OF RIGHT EPIDIDYMIS|MALIGNANT NEOPLASM OF RIGHT EPIDIDYMIS
C2845881|T191|C63.00|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED EPIDIDYMIS|MALIGNANT NEOPLASM OF UNSPECIFIED EPIDIDYMIS
C2861588|T191|C92.22|ICD10CM|ATYPICAL CHRONIC MYELOID LEUKEMIA, BCR/ABL-NEGATIVE, IN RELAPSE|ATYPICAL CHRONIC MYELOID LEUKEMIA, BCR/ABL-NEG, IN RELAPSE
C2905709|T037|X74.09XS|ICD10CM|INTENTIONAL SELF-HARM BY OTHER GAS, AIR OR SPRING-OPERATED GUN, SEQUELA|SELF-HARM BY OTH GAS, AIR OR SPRING-OPERATED GUN, SEQUELA
C2875026|T047|G04.91|ICD10CM|MYELITIS, UNSPECIFIED|MYELITIS, UNSPECIFIED
C2905708|T037|X74.09XD|ICD10CM|INTENTIONAL SELF-HARM BY OTHER GAS, AIR OR SPRING-OPERATED GUN, SUBSEQUENT ENCOUNTER|SELF-HARM BY OTH GAS, AIR OR SPRING-OPERATED GUN, SUBS
C4268033|T047|E10.3493|ICD10CM|TYPE 1 DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|TYPE 1 DIAB WITH SEVERE NONP RTNOP WITHOUT MACULAR EDEMA, BI
C2887936|T047|K72.90|ICD10CM|HEPATIC FAILURE, UNSPECIFIED WITHOUT COMA|HEPATIC FAILURE, UNSPECIFIED WITHOUT COMA
C4268031|T047|E10.3491|ICD10CM|TYPE 1 DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|TYPE 1 DIAB WITH SEVERE NONP RTNOP WITHOUT MCLR EDEMA, R EYE
C2853902|T191||ICD10CM|MANTLE CELL LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES
C2890863|T037|T84.621A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL FIXATION DEVICE OF LEFT FEMUR, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INT FIX OF LEFT FEMUR, INIT
C4268034|T047|E10.3499|ICD10CM|TYPE 1 DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|TYPE 1 DIAB WITH SEVERE NONP RTNOP WITHOUT MCLR EDEMA, UNSP
C4270447|T046|T83.86XA|ICD10CM|THROMBOSIS DUE TO GENITOURINARY PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|THROMBOSIS DUE TO GENITOURINARY PROSTH DEV/GRFT, INIT
C2874575|T048||ICD10CM|COCAINE ABUSE WITH INTOXICATION, UNCOMPLICATED
C2879233|T037|T45.612S|ICD10CM|POISONING BY THROMBOLYTIC DRUG, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY THROMBOLYTIC DRUG, SELF-HARM, SEQUELA
C2874424|T048|F11.121|ICD10CM|OPIOID ABUSE WITH INTOXICATION DELIRIUM|OPIOID ABUSE WITH INTOXICATION DELIRIUM
C2858234|T037|S72.391A|ICD10CM|OTHER FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF SHAFT OF RIGHT FEMUR, INIT FOR CLOS FX
C4267998|T047|E09.3551|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, RIGHT EYE|DRUG/CHEM DIABETES WITH STABLE PROLIF DIABETIC RTNOP, R EYE
C4267999|T047|E09.3552|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, LEFT EYE|DRUG/CHEM DIAB WITH STABLE PROLIF DIABETIC RTNOP, LEFT EYE
C4268000|T047|E09.3553|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, BILATERAL|DRUG/CHEM DIABETES WITH STABLE PROLIF DIABETIC RTNOP, BI
C2832453|T037|S06.4X6A|ICD10CM|EPIDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|EPIDURAL HEMORRHAGE W LOC >24 HR W/O RET CONSC W SURV, INIT
C4268001|T047|E09.3559|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, UNSPECIFIED EYE|DRUG/CHEM DIABETES WITH STABLE PROLIF DIABETIC RTNOP, UNSP
C2879231|T037|T45.612A|ICD10CM|POISONING BY THROMBOLYTIC DRUG, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY THROMBOLYTIC DRUG, INTENTIONAL SELF-HARM, INIT
C2876619|T037|T36.3X2A|ICD10CM|POISONING BY MACROLIDES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY MACROLIDES, INTENTIONAL SELF-HARM, INIT ENCNTR
C2835290|T037|S22.039A|ICD10CM|UNSPECIFIED FRACTURE OF THIRD THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF THIRD THORACIC VERTEBRA, INIT FOR CLOS FX
C2835291|T037|S22.039B|ICD10CM|UNSPECIFIED FRACTURE OF THIRD THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF THIRD THORACIC VERTEBRA, INIT FOR OPN FX
C2902160|T046|M87.869|ICD10CM|OTHER OSTEONECROSIS, UNSPECIFIED FIBULA|OTHER OSTEONECROSIS, UNSPECIFIED FIBULA
C2902156|T046|M87.862|ICD10CM|OTHER OSTEONECROSIS, LEFT TIBIA|OTHER OSTEONECROSIS, LEFT TIBIA
C2902157|T046|M87.863|ICD10CM|OTHER OSTEONECROSIS, UNSPECIFIED TIBIA|OTHER OSTEONECROSIS, UNSPECIFIED TIBIA
C2902155|T046|M87.861|ICD10CM|OTHER OSTEONECROSIS, RIGHT TIBIA|OTHER OSTEONECROSIS, RIGHT TIBIA
C2896589|T046|M80.059A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, UNSP FEMUR, INIT
C2902158|T046|M87.864|ICD10CM|OTHER OSTEONECROSIS, RIGHT FIBULA|OTHER OSTEONECROSIS, RIGHT FIBULA
C2902159|T046|M87.865|ICD10CM|OTHER OSTEONECROSIS, LEFT FIBULA|OTHER OSTEONECROSIS, LEFT FIBULA
C2832022|T037|S06.2X2S|ICD10CM|DIFFUSE TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|DIFFUSE TBI W LOSS OF CONSCIOUSNESS OF 31-59 MIN, SEQUELA
C2886741|T037|T79.7XXA|ICD10CM|TRAUMATIC SUBCUTANEOUS EMPHYSEMA, INITIAL ENCOUNTER|TRAUMATIC SUBCUTANEOUS EMPHYSEMA, INITIAL ENCOUNTER
C0348589|T047|I23.8|DMDICD10|OTHER CURRENT COMPLICATIONS FOLLOWING ACUTE MYOCARDIAL INFARCTION|SONSTIGE AKUTE KOMPLIKATIONEN NACH AKUTEM MYOKARDINFARKT
C2874856|T048|F19.99|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH UNSPECIFIED PSYCHOACTIVE SUBSTANCE-INDUCED DISORDER|OTH PSYCHOACTIVE SUBSTANCE USE, UNSP W UNSP DISORDER
C2874850|T048|F19.96|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH PSYCHOACTIVE SUBSTANCE-INDUCED PERSISTING AMNESTIC DISORDER|OTH PSYCHOACTV SUB USE, UNSP W PERSIST AMNESTIC DISORDER
C4237273|T048|F19.97|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH PSYCHOACTIVE SUBSTANCE-INDUCED PERSISTING DEMENTIA|OTHER (OR UNKNOWN) SUBSTANCE-INDUCED MAJOR NEUROCOGNITIVE DISORDER, WITHOUT USE DISORDER
C4268299|T048|F19.94|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH PSYCHOACTIVE SUBSTANCE-INDUCED MOOD DISORDER|OTHER (OR UNKNOWN) SUBSTANCE-INDUCED BIPOLAR OR RELATED DISORDER, WITHOUT USE DISORDER
C1142492|T046|I23.7|ICD10CM|POSTINFARCTION ANGINA|POSTINFARCTION ANGINA
C0348865|T046|I23.0|DMDICD10|HEMOPERICARDIUM AS CURRENT COMPLICATION FOLLOWING ACUTE MYOCARDIAL INFARCTION|HAEMOPERIKARD ALS AKUTE KOMPLIKATION NACH AKUTEM MYOKARDINFARKT
C0348866|T047|I23.1|DMDICD10|ATRIAL SEPTAL DEFECT AS CURRENT COMPLICATION FOLLOWING ACUTE MYOCARDIAL INFARCTION|VORHOFSEPTUMDEFEKT ALS AKUTE KOMPLIKATION NACH AKUTEM MYOKARDINFARKT
C0340331|T047|I23.2|DMDICD10|VENTRICULAR SEPTAL DEFECT AS CURRENT COMPLICATION FOLLOWING ACUTE MYOCARDIAL INFARCTION|VENTRIKELSEPTUMDEFEKT ALS AKUTE KOMPLIKATION NACH AKUTEM MYOKARDINFARKT
C0348867|T047|I23.3|DMDICD10|RUPTURE OF CARDIAC WALL WITHOUT HEMOPERICARDIUM AS CURRENT COMPLICATION FOLLOWING ACUTE MYOCARDIAL INFARCTION|RUPTUR DER HERZWAND OHNE HAEMOPERIKARD ALS AKUTE KOMPLIKATION NACH AKUTEM MYOKARDINFARKT
C2832020|T037|S06.2X2A|ICD10CM|DIFFUSE TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|DIFFUSE TBI W LOSS OF CONSCIOUSNESS OF 31-59 MIN, INIT
C2890406|T037|T84.011A|ICD10CM|BROKEN INTERNAL LEFT HIP PROSTHESIS, INITIAL ENCOUNTER|BROKEN INTERNAL LEFT HIP PROSTHESIS, INITIAL ENCOUNTER
C2833502|T037|S12.490A|ICD10CM|OTHER DISPLACED FRACTURE OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH DISP FX OF FIFTH CERVICAL VERTEBRA, INIT FOR CLOS FX
C2833503|T037|S12.490B|ICD10CM|OTHER DISPLACED FRACTURE OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH DISP FX OF FIFTH CERVICAL VERTEBRA, INIT FOR OPN FX
C2858961|T037|S72.472A|ICD10CM|TORUS FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TORUS FRACTURE OF LOWER END OF LEFT FEMUR, INIT FOR CLOS FX
C0477745|T047|N17.8|DMDICD10|OTHER ACUTE KIDNEY FAILURE|SONSTIGES AKUTES NIERENVERSAGEN
C2890115|T037|T82.594A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INFUSION CATHETER, INITIAL ENCOUNTER|MECH COMPL OF INFUSION CATHETER, INITIAL ENCOUNTER
C2874487|T048|F12.222|ICD10CM|CANNABIS DEPENDENCE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE|CANNABIS DEPENDENCE W INTOXICATION W PERCEPTUAL DISTURBANCE
C2874486|T048|F12.221|ICD10CM|CANNABIS DEPENDENCE WITH INTOXICATION DELIRIUM|CANNABIS DEPENDENCE WITH INTOXICATION DELIRIUM
C2874485|T048||ICD10CM|CANNABIS DEPENDENCE WITH INTOXICATION, UNCOMPLICATED
C2832649|T037|S06.894S|ICD10CM|OTHER SPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|INTCRAN INJ W LOC OF 6 HOURS TO 24 HOURS, SEQUELA
C2889395|T047|M06.032|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, LEFT WRIST|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, LEFT WRIST
C2874488|T048|F12.229|ICD10CM|CANNABIS DEPENDENCE WITH INTOXICATION, UNSPECIFIED|CANNABIS DEPENDENCE WITH INTOXICATION, UNSPECIFIED
C2889394|T047|M06.031|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, RIGHT WRIST|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, RIGHT WRIST
C2857927|T037|S72.341C|ICD10CM|DISPLACED SPIRAL FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL SPIRAL FX SHAFT OF R FEMR, INIT FOR OPN FX TYPE 3A/B/C
C2832016|T037|S06.2X1A|ICD10CM|DIFFUSE TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|DIFFUSE TBI W LOC OF 30 MINUTES OR LESS, INIT
C2885061|T037|T60.3X2S|ICD10CM|TOXIC EFFECT OF HERBICIDES AND FUNGICIDES, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF HERBICIDES AND FUNGICIDES, SLF-HRM, SEQUELA
C2832401|T037|S06.383S|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF BRAINSTEM WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, SEQUELA|CONTUS/LAC/HEM BRAINSTEM W LOC OF 1-5 HRS 59 MIN, SEQUELA
C2832272|T037|S06.352S|ICD10CM|TRAUMATIC HEMORRHAGE OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|TRAUM HEMOR LEFT CEREBRUM W LOC OF 31-59 MIN, SEQUELA
C2855851|T037|S68.021S|ICD10CM|PARTIAL TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF RIGHT THUMB, SEQUELA|PARTIAL TRAUMATIC MCP AMPUTATION OF RIGHT THUMB, SEQUELA
C2838606|T037|S34.01XD|ICD10CM|CONCUSSION AND EDEMA OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|CONCUSSION AND EDEMA OF LUMBAR SPINAL CORD, SUBS ENCNTR
C4269497|T037|S02.632B|ICD10CM|FRACTURE OF CORONOID PROCESS OF LEFT MANDIBLE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF CORONOID PROCESS OF LEFT MANDIBLE, 7THB
C2832270|T037|S06.352A|ICD10CM|TRAUMATIC HEMORRHAGE OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|TRAUM HEMOR LEFT CEREBRUM W LOC OF 31-59 MIN, INIT
C2837897|T037|S32.402A|ICD10CM|UNSPECIFIED FRACTURE OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF LEFT ACETABULUM, INIT FOR CLOS FX
C2837898|T037|S32.402B|ICD10CM|UNSPECIFIED FRACTURE OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF LEFT ACETABULUM, INIT FOR OPN FX
C2890475|T037|T84.039A|ICD10CM|MECHANICAL LOOSENING OF UNSPECIFIED INTERNAL PROSTHETIC JOINT, INITIAL ENCOUNTER|MECHANICAL LOOSENING OF UNSP INTERNAL PROSTHETIC JOINT, INIT
C4270239|T046|T83.092A|ICD10CM|OTHER MECHANICAL COMPLICATION OF NEPHROSTOMY CATHETER, INITIAL ENCOUNTER|MECH COMPL OF NEPHROSTOMY CATHETER, INITIAL ENCOUNTER
C2901819|T047|M86.219|ICD10CM|SUBACUTE OSTEOMYELITIS, UNSPECIFIED SHOULDER|SUBACUTE OSTEOMYELITIS, UNSPECIFIED SHOULDER
C2878382|T037|T43.212S|ICD10CM|POISONING BY SELECTIVE SEROTONIN AND NOREPINEPHRINE REUPTAKE INHIBITORS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY SLCTV SEROTON/NOREPINEPH REUP INHIBTR,SLF-HRM, SQLA
C2901821|T047|M86.212|ICD10CM|SUBACUTE OSTEOMYELITIS, LEFT SHOULDER|SUBACUTE OSTEOMYELITIS, LEFT SHOULDER
C2901820|T047|M86.211|ICD10CM|SUBACUTE OSTEOMYELITIS, RIGHT SHOULDER|SUBACUTE OSTEOMYELITIS, RIGHT SHOULDER
C2869844|T037|S98.219S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF TWO OR MORE UNSPECIFIED LESSER TOES, SEQUELA|COMPLETE TRAUM AMP OF TWO OR MORE UNSP LESSER TOES, SEQUELA
C2882378|T047|I63.349|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF UNSPECIFIED CEREBELLAR ARTERY|CEREBRAL INFARCTION DUE TO THOMBOS UNSP CEREBELLAR ARTERY
C2878380|T037|T43.212A|ICD10CM|POISONING BY SELECTIVE SEROTONIN AND NOREPINEPHRINE REUPTAKE INHIBITORS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY SLCTV SEROTON/NOREPINEPH REUP INHIBTR,SLF-HRM, INIT
C2882376|T047|I63.341|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF RIGHT CEREBELLAR ARTERY|CEREBRAL INFRC DUE TO THROMBOSIS OF RIGHT CEREBLR ARTERY
C4268484|T047|I63.343|ICD10CM|CEREBRAL INFARCTION TO THROMBOSIS OF BILATERAL CEREBELLAR ARTERIES|CEREBRAL INFRC TO THROMBOSIS OF BILATERAL CEREBLR ARTERIES
C2882377|T047|I63.342|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF LEFT CEREBELLAR ARTERY|CEREBRAL INFARCTION DUE TO THROMBOSIS OF LEFT CEREBLR ARTERY
C2884054|T037|T51.8X2S|ICD10CM|TOXIC EFFECT OF OTHER ALCOHOLS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF OTH ALCOHOLS, INTENTIONAL SELF-HARM, SEQUELA
C2861582|T191|C92.10|ICD10CM|CHRONIC MYELOID LEUKEMIA, BCR/ABL-POSITIVE, NOT HAVING ACHIEVED REMISSION|CHRONIC MYELOID LEUK, BCR/ABL-POSITIVE, NOT ACHIEVE REMIS
C2861583|T191|C92.11|ICD10CM|CHRONIC MYELOID LEUKEMIA, BCR/ABL-POSITIVE, IN REMISSION|CHRONIC MYELOID LEUKEMIA, BCR/ABL-POSITIVE, IN REMISSION
C2861584|T191|C92.12|ICD10CM|CHRONIC MYELOID LEUKEMIA, BCR/ABL-POSITIVE, IN RELAPSE|CHRONIC MYELOID LEUKEMIA, BCR/ABL-POSITIVE, IN RELAPSE
C0837606|T046|M06.39|ICD10AM|RHEUMATOID NODULE, MULTIPLE SITES|RHEUMATOID NODULE, SITE UNSPECIFIED
C2889465|T046|M06.38|ICD10CM|RHEUMATOID NODULE, VERTEBRAE|RHEUMATOID NODULE, VERTEBRAE
C2876768|T037|T36.92XA|ICD10CM|POISONING BY UNSPECIFIED SYSTEMIC ANTIBIOTIC, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY UNSP SYSTEMIC ANTIBIOTIC, SELF-HARM, INIT
C0837606|T046||ICD10CM|RHEUMATOID NODULE, UNSPECIFIED SITE
C2833999|T037|S14.142S|ICD10CM|BROWN-SEQUARD SYNDROME AT C2 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|BROWN-SEQUARD SYNDROME AT C2, SEQUELA
C2856932|T037|S72.059C|ICD10CM|UNSPECIFIED FRACTURE OF HEAD OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP FX HEAD OF UNSP FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2856931|T037|S72.059B|ICD10CM|UNSPECIFIED FRACTURE OF HEAD OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP FX HEAD OF UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C4268233|T048|F14.14|ICD10CM|COCAINE ABUSE WITH COCAINE-INDUCED MOOD DISORDER|COCAINE USE DISORDER, MILD, WITH COCAINE-INDUCED DEPRESSIVE DISORDER
C2889647|T047|M08.962|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, LEFT KNEE|JUVENILE ARTHRITIS, UNSPECIFIED, LEFT KNEE
C2895359|T047|M49.88|ICD10CM|SPONDYLOPATHY IN DISEASES CLASSIFIED ELSEWHERE, SACRAL AND SACROCOCCYGEAL REGION|SPOND IN DISEASES CLASSD ELSWHR, SACR/SACROCYGL REGION
C2889646|T047|M08.961|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, RIGHT KNEE|JUVENILE ARTHRITIS, UNSPECIFIED, RIGHT KNEE
C0494735|T047|K28.6|DMDICD10|CHRONIC OR UNSPECIFIED GASTROJEJUNAL ULCER WITH BOTH HEMORRHAGE AND PERFORATION|ULCUS PEPTICUM JEJUNI: CHRONISCH ODER NICHT NAEHER BEZEICHNET, MIT BLUTUNG UND PERFORATION
C2889648|T047|M08.969|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, UNSPECIFIED KNEE|JUVENILE ARTHRITIS, UNSPECIFIED, UNSPECIFIED KNEE
C4270368|T046|T83.711A|ICD10CM|EROSION OF IMPLANTED VAGINAL MESH TO SURROUNDING ORGAN OR TISSUE, INITIAL ENCOUNTER|EROSN IMPLNT VAGINAL MESH TO SURRND ORG/TISS, INIT
C2858355|T037|S72.412A|ICD10CM|DISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED UNSP CONDYLE FX LOWER END OF LEFT FEMUR, INIT
C2858356|T037|S72.412B|ICD10CM|DISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL UNSP CONDYLE FX LOW END L FEMR, 7THB
C2858357|T037|S72.412C|ICD10CM|DISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL UNSP CONDYLE FX LOW END L FEMR, 7THC
C4268394|T047|H35.3293|ICD10CM|EXUDATIVE AGE-RELATED MACULAR DEGENERATION, UNSPECIFIED EYE, WITH INACTIVE SCAR|EXUDATIVE AGE-RELATED MCLR DEGN, UNSP, WITH INACTIVE SCAR
C4268393|T047|H35.3292|ICD10CM|EXUDATIVE AGE-RELATED MACULAR DEGENERATION, UNSPECIFIED EYE, WITH INACTIVE CHOROIDAL NEOVASCULARIZATION|EXUDATIVE AGE-REL MCLR DEGN, UNSP, WITH INACT CHRDL NEOVAS
C4268392|T047|H35.3291|ICD10CM|EXUDATIVE AGE-RELATED MACULAR DEGENERATION, UNSPECIFIED EYE, WITH ACTIVE CHOROIDAL NEOVASCULARIZATION|EXUDATIVE AGE-REL MCLR DEGN, UNSP, WITH ACTV CHRDL NEOVAS
C4268391|T047|H35.3290|ICD10CM|EXUDATIVE AGE-RELATED MACULAR DEGENERATION, UNSPECIFIED EYE, STAGE UNSPECIFIED|EXUDATIVE AGE-RELATED MCLR DEGN, UNSP, STAGE UNSPECIFIED
C0007115|T191|C73|DMDICD10|MALIGNANT NEOPLASM OF THYROID GLAND|BOESARTIGE NEUBILDUNG DER SCHILDDRUESE
C4268107|T047|E11.3541|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, RIGHT EYE|TYPE 2 DIAB WITH PROLIF DIAB RTNOP WITH COMB DETACH, R EYE
C4268108|T047|E11.3542|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, LEFT EYE|TYPE 2 DIAB WITH PROLIF DIAB RTNOP WITH COMB DETACH, L EYE
C4268109|T047|E11.3543|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, BILATERAL|TYPE 2 DIAB WITH PROLIF DIABETIC RTNOP WITH COMB DETACH, BI
C2888653|T047|L97.123|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT THIGH WITH NECROSIS OF MUSCLE|NON-PRS CHRONIC ULCER OF LEFT THIGH W NECROSIS OF MUSCLE
C4268110|T047|E11.3549|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, UNSPECIFIED EYE|TYPE 2 DIAB WITH PROLIF DIAB RTNOP WITH COMB DETACH, UNSP
C2831996|T037|S06.1X6A|ICD10CM|TRAUMATIC CEREBRAL EDEMA WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|TRAUM CEREBRAL EDEMA W LOC >24 HR W/O RET CONSC W SURV, INIT
C2910838|T033|Z44.101|ICD10CM|ENCOUNTER FOR FITTING AND ADJUSTMENT OF UNSPECIFIED RIGHT ARTIFICIAL LEG|ENCOUNTER FOR FIT/ADJST OF UNSP RIGHT ARTIFICIAL LEG
C2910839|T033|Z44.102|ICD10CM|ENCOUNTER FOR FITTING AND ADJUSTMENT OF UNSPECIFIED LEFT ARTIFICIAL LEG|ENCOUNTER FOR FIT/ADJST OF UNSP LEFT ARTIFICIAL LEG
C2910840|T033|Z44.109|ICD10CM|ENCOUNTER FOR FITTING AND ADJUSTMENT OF UNSPECIFIED ARTIFICIAL LEG, UNSPECIFIED LEG|ENCOUNTER FOR FIT/ADJST OF UNSP ARTIFICIAL LEG, UNSP LEG
C2831998|T037|S06.1X6S|ICD10CM|TRAUMATIC CEREBRAL EDEMA WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|TRAUM CEREB EDEMA W LOC >24 HR W/O RET CONSC W SURV, SEQUELA
C0020255|T047|G91.9|DMDICD10|HYDROCEPHALUS, UNSPECIFIED|HYDROZEPHALUS, NICHT NAEHER BEZEICHNET
C0477417|T047|G91.8|DMDICD10|OTHER HYDROCEPHALUS|SONSTIGER HYDROZEPHALUS
C2886771|T037|T79.A3XA|ICD10CM|TRAUMATIC COMPARTMENT SYNDROME OF ABDOMEN, INITIAL ENCOUNTER|TRAUMATIC COMPARTMENT SYNDROME OF ABDOMEN, INITIAL ENCOUNTER
C0477432|T047|G91.3|DMDICD10|POST-TRAUMATIC HYDROCEPHALUS, UNSPECIFIED|POSTTRAUMATISCHER HYDROZEPHALUS, NICHT NAEHER BEZEICHNET
C2047886|T047||ICD10CM|(IDIOPATHIC) NORMAL PRESSURE HYDROCEPHALUS
C0549423|T047|G91.1|DMDICD10|OBSTRUCTIVE HYDROCEPHALUS|HYDROCEPHALUS OCCLUSUS
C1955759|T047||ICD10CM|COMMUNICATING HYDROCEPHALUS
C2833890|T037|S14.113A|ICD10CM|COMPLETE LESION AT C3 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION AT C3 LEVEL OF CERVICAL SPINAL CORD, INIT
C2859186|T037|S73.021A|ICD10CM|OBTURATOR SUBLUXATION OF RIGHT HIP, INITIAL ENCOUNTER|OBTURATOR SUBLUXATION OF RIGHT HIP, INITIAL ENCOUNTER
C2875379|T047|G91.4|ICD10CM|HYDROCEPHALUS IN DISEASES CLASSIFIED ELSEWHERE|HYDROCEPHALUS IN DISEASES CLASSIFIED ELSEWHERE
C2832692|T037|S06.9X5A|ICD10CM|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, INITIAL ENCOUNTER|UNSP INTRACRANIAL INJURY W LOC >24 HR W RET CONSC LEV, INIT
C2895356|T047|M49.85|ICD10CM|SPONDYLOPATHY IN DISEASES CLASSIFIED ELSEWHERE, THORACOLUMBAR REGION|SPOND IN DISEASES CLASSD ELSWHR, THORACOLUMBAR REGION
C2833892|T037|S14.113S|ICD10CM|COMPLETE LESION AT C3 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|COMPLETE LESION AT C3 LEVEL OF CERVICAL SPINAL CORD, SEQUELA
C2843299|T037|S48.112A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN LEFT SHOULDER AND ELBOW, INITIAL ENCOUNTER|COMPLETE TRAUM AMP AT LEVEL BETW L SHOULDER AND ELBOW, INIT
C4269208|T033|R40.2432|ICD10CM|GLASGOW COMA SCALE SCORE 3-8, AT ARRIVAL TO EMERGENCY DEPARTMENT|GLASGOW COMA SCALE SCORE 3-8, EMR
C4269209|T033|R40.2433|ICD10CM|GLASGOW COMA SCALE SCORE 3-8, AT HOSPITAL ADMISSION|GLASGOW COMA SCALE SCORE 3-8, AT HOSPITAL ADMISSION
C4269206|T033|R40.2430|ICD10CM|GLASGOW COMA SCALE SCORE 3-8, UNSPECIFIED TIME|GLASGOW COMA SCALE SCORE 3-8, UNSPECIFIED TIME
C4269207|T033|R40.2431|ICD10CM|GLASGOW COMA SCALE SCORE 3-8, IN THE FIELD [EMT OR AMBULANCE]|GLASGOW COMA SCALE SCORE 3-8, IN THE FIELD
C2905726|T037|X77.0XXA|ICD10CM|INTENTIONAL SELF-HARM BY STEAM OR HOT VAPORS, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY STEAM OR HOT VAPORS, INIT ENCNTR
C2878173|T037|T42.5X2A|ICD10CM|POISONING BY MIXED ANTIEPILEPTICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY MIXED ANTIEPILEPTICS, SELF-HARM, INIT
C4269210|T033|R40.2434|ICD10CM|GLASGOW COMA SCALE SCORE 3-8, 24 HOURS OR MORE AFTER HOSPITAL ADMISSION|GLASGOW COMA SCALE SCORE 3-8, 24+HRS
C2865574|T037|S88.912S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT LOWER LEG, LEVEL UNSPECIFIED, SEQUELA|COMPLETE TRAUMATIC AMP OF L LOW LEG, LEVEL UNSP, SEQUELA
C2890742|T037|T84.298A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTERNAL FIXATION DEVICE OF OTHER BONES, INITIAL ENCOUNTER|MECH COMPL OF INTERNAL FIXATION DEVICE OF OTH BONES, INIT
C2843301|T037|S48.112S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN LEFT SHOULDER AND ELBOW, SEQUELA|COMPLETE TRAUM AMP AT LEVEL BETW L SHLDR AND ELBOW, SEQUELA
C2835154|T037|S22.000A|ICD10CM|WEDGE COMPRESSION FRACTURE OF UNSPECIFIED THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|WEDGE COMPRESSION FRACTURE OF UNSP THORACIC VERTEBRA, INIT
C2835155|T037|S22.000B|ICD10CM|WEDGE COMPRESSION FRACTURE OF UNSPECIFIED THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|WEDGE COMPRSN FX UNSP THOR VERTEBRA, INIT FOR OPN FX
C2835847|T037|S24.152S|ICD10CM|OTHER INCOMPLETE LESION AT T2-T6 LEVEL OF THORACIC SPINAL CORD, SEQUELA|OTH INCOMPLETE LESION AT T2-T6, SEQUELA
C2865573|T037|S88.912D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT LOWER LEG, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF L LOW LEG, LEVEL UNSP, SUBS
C2895355|T047|M49.84|ICD10CM|SPONDYLOPATHY IN DISEASES CLASSIFIED ELSEWHERE, THORACIC REGION|SPONDYLOPATHY IN DISEASES CLASSD ELSWHR, THORACIC REGION
C2865572|T037|S88.912A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT LOWER LEG, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF L LOW LEG, LEVEL UNSP, INIT
C2905728|T037|X77.0XXS|ICD10CM|INTENTIONAL SELF-HARM BY STEAM OR HOT VAPORS, SEQUELA|INTENTIONAL SELF-HARM BY STEAM OR HOT VAPORS, SEQUELA
C2878175|T037|T42.5X2S|ICD10CM|POISONING BY MIXED ANTIEPILEPTICS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY MIXED ANTIEPILEPTICS, SELF-HARM, SEQUELA
C2835784|T037|S24.113A|ICD10CM|COMPLETE LESION AT T7-T10 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION AT T7-T10, INIT
C2835785|T037|S24.113D|ICD10CM|COMPLETE LESION AT T7-T10 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION AT T7-T10, SUBS
C2883836|T037|T50.A22A|ICD10CM|POISONING BY MIXED BACTERIAL VACCINES WITHOUT A PERTUSSIS COMPONENT, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY MIXED BACT VACCINES W/O A PERTUSS, SELF-HARM, INIT
C4268948|T046|N99.521|ICD10CM|INFECTION OF INCONTINENT EXTERNAL STOMA OF URINARY TRACT|INFECTION OF INCONTINENT EXTERNAL STOMA OF URINARY TRACT
C4268947|T046|N99.520|ICD10CM|HEMORRHAGE OF INCONTINENT EXTERNAL STOMA OF URINARY TRACT|HEMORRHAGE OF INCONTINENT EXTERNAL STOMA OF URINARY TRACT
C4268950|T046|N99.523|ICD10CM|HERNIATION OF INCONTINENT STOMA OF URINARY TRACT|HERNIATION OF INCONTINENT STOMA OF URINARY TRACT
C4268949|T046|N99.522|ICD10CM|MALFUNCTION OF INCONTINENT EXTERNAL STOMA OF URINARY TRACT|MALFUNCTION OF INCONTINENT EXTERNAL STOMA OF URINARY TRACT
C4268951|T046|N99.524|ICD10CM|STENOSIS OF INCONTINENT STOMA OF URINARY TRACT|STENOSIS OF INCONTINENT STOMA OF URINARY TRACT
C2883838|T037|T50.A22S|ICD10CM|POISONING BY MIXED BACTERIAL VACCINES WITHOUT A PERTUSSIS COMPONENT, INTENTIONAL SELF-HARM, SEQUELA|POISN BY MIXED BACT VACCINES W/O A PERTUSS, SLF-HRM, SEQUELA
C4268952|T046|N99.528|ICD10CM|OTHER COMPLICATION OF INCONTINENT EXTERNAL STOMA OF URINARY TRACT|OTHER COMP OF INCONTINENT EXTERNAL STOMA OF URINARY TRACT
C2882699|T047|I70.213|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES WITH INTERMITTENT CLAUDICATION, BILATERAL LEGS|ATHSCL NATIVE ARTERIES OF EXTRM W INTRMT CLAUD, BI LEGS
C2882698|T047|I70.212|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES WITH INTERMITTENT CLAUDICATION, LEFT LEG|ATHSCL NATIVE ARTERIES OF EXTRM W INTRMT CLAUD, LEFT LEG
C2882697|T047|I70.211|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES WITH INTERMITTENT CLAUDICATION, RIGHT LEG|ATHSCL NATIVE ARTERIES OF EXTRM W INTRMT CLAUD, RIGHT LEG
C2889140|T047|M05.122|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT ELBOW|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2890706|T037|T84.218A|ICD10CM|BREAKDOWN (MECHANICAL) OF INTERNAL FIXATION DEVICE OF OTHER BONES, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF INT FIX OF BONES, INIT
C2889141|T047|M05.129|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP ELBOW
C2882701|T047|I70.219|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES WITH INTERMITTENT CLAUDICATION, UNSPECIFIED EXTREMITY|ATHSCL NATIVE ARTERIES OF EXTRM W INTRMT CLAUD, UNSP EXTRM
C2882700|T047|I70.218|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES WITH INTERMITTENT CLAUDICATION, OTHER EXTREMITY|ATHSCL NATIVE ARTERIES OF EXTRM W INTRMT CLAUD, OTH EXTRM
C2874068|T047||ICD10CM|TYPE 1 DIABETES MELLITUS WITH HYPOGLYCEMIA WITH COMA
C2888621|T047|L89.91|ICD10CM|PRESSURE ULCER OF UNSPECIFIED SITE, STAGE 1|PRESSURE ULCER OF UNSPECIFIED SITE, STAGE 1
C2874069|T047||ICD10CM|TYPE 1 DIABETES MELLITUS WITH HYPOGLYCEMIA WITHOUT COMA
C2901452|T046|M84.641A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, RIGHT HAND, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, RIGHT HAND, INIT
C2874440|T048|F11.222|ICD10CM|OPIOID DEPENDENCE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE|OPIOID DEPENDENCE W INTOXICATION WITH PERCEPTUAL DISTURBANCE
C2837825|T037|S32.311A|ICD10CM|DISPLACED AVULSION FRACTURE OF RIGHT ILIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED AVULSION FRACTURE OF RIGHT ILIUM, INIT FOR CLOS FX
C2874438|T048||ICD10CM|OPIOID DEPENDENCE WITH INTOXICATION, UNCOMPLICATED
C2874439|T048|F11.221|ICD10CM|OPIOID DEPENDENCE WITH INTOXICATION DELIRIUM|OPIOID DEPENDENCE WITH INTOXICATION DELIRIUM
C2884122|T037|T52.2X2S|ICD10CM|TOXIC EFFECT OF HOMOLOGUES OF BENZENE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF HOMOLOGUES OF BENZENE, SELF-HARM, SEQUELA
C2884102|T037|T52.1X2A|ICD10CM|TOXIC EFFECT OF BENZENE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF BENZENE, INTENTIONAL SELF-HARM, INIT ENCNTR
C2874441|T048|F11.229|ICD10CM|OPIOID DEPENDENCE WITH INTOXICATION, UNSPECIFIED|OPIOID DEPENDENCE WITH INTOXICATION, UNSPECIFIED
C4269343|T037|S02.31XB|ICD10CM|FRACTURE OF ORBITAL FLOOR, RIGHT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF ORBITAL FLOOR, RIGHT SIDE, 7THB
C4269342|T037|S02.31XA|ICD10CM|FRACTURE OF ORBITAL FLOOR, RIGHT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF ORBITAL FLOOR, RIGHT SIDE, INIT
C2886366|T037|T71.132S|ICD10CM|ASPHYXIATION DUE TO BEING TRAPPED IN BED LINENS, INTENTIONAL SELF-HARM, SEQUELA|ASPHYX DUE TO BEING TRAPPED IN BED LINENS, SLF-HRM, SEQUELA
C2890254|T037|T83.118A|ICD10CM|BREAKDOWN (MECHANICAL) OF OTHER URINARY DEVICES AND IMPLANTS, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF URINARY DEVICES AND IMPLANTS, INIT
C2884104|T037|T52.1X2S|ICD10CM|TOXIC EFFECT OF BENZENE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF BENZENE, INTENTIONAL SELF-HARM, SEQUELA
C2884120|T037|T52.2X2A|ICD10CM|TOXIC EFFECT OF HOMOLOGUES OF BENZENE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF HOMOLOGUES OF BENZENE, SELF-HARM, INIT
C4269347|T037|S02.31XS|ICD10CM|FRACTURE OF ORBITAL FLOOR, RIGHT SIDE, SEQUELA|FRACTURE OF ORBITAL FLOOR, RIGHT SIDE, SEQUELA
C2860031|T037|S78.919A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED HIP AND THIGH, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|COMPLETE TRAUM AMP OF UNSP HIP AND THIGH, LEVEL UNSP, INIT
C2860032|T037|S78.919D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED HIP AND THIGH, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|COMPLETE TRAUM AMP OF UNSP HIP AND THIGH, LEVEL UNSP, SUBS
C2860033|T037|S78.919S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED HIP AND THIGH, LEVEL UNSPECIFIED, SEQUELA|COMPLETE TRAUM AMP OF UNSP HIP AND THIGH, LEVEL UNSP, SQLA
C2833197|T037|S12.090A|ICD10CM|OTHER DISPLACED FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH DISP FX OF FIRST CERVICAL VERTEBRA, INIT FOR CLOS FX
C2833198|T037|S12.090B|ICD10CM|OTHER DISPLACED FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH DISP FX OF FIRST CERVICAL VERTEBRA, INIT FOR OPN FX
C0868576|T033||ICD10CM|OTHER ARTIFICIAL OPENINGS OF URINARY TRACT STATUS
C2977944|T191|C72.9|ICD10CM|MALIGNANT NEOPLASM OF CENTRAL NERVOUS SYSTEM, UNSPECIFIED|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF CENTRAL NERVOUS SYSTEM
C0496760|T191|C05.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF PALATE|BOESARTIGE NEUBILDUNG: GAUMEN, MEHRERE TEILBEREICHE UEBERLAPPEND
C0153378|T191|C05.9|DMDICD10|MALIGNANT NEOPLASM OF PALATE, UNSPECIFIED|BOESARTIGE NEUBILDUNG: GAUMEN, NICHT NAEHER BEZEICHNET
C0153646|T191|C72.0|DMDICD10|MALIGNANT NEOPLASM OF SPINAL CORD|BOESARTIGE NEUBILDUNG: RUECKENMARK
C0349017|T191|C72.1|DMDICD10|MALIGNANT NEOPLASM OF CAUDA EQUINA|BOESARTIGE NEUBILDUNG: CAUDA EQUINA
C2521566|T060|C050|ICD10PCS|MALIGNANT NEOPLASM OF HARD PALATE|NUCLEAR MEDICINE @ CENTRAL NERVOUS SYSTEM @ NONIMAGING NUCLEAR MEDICINE PROBE @ BRAIN
C0153376|T191|C05.1|DMDICD10|MALIGNANT NEOPLASM OF SOFT PALATE|BOESARTIGE NEUBILDUNG: WEICHER GAUMEN
C4509292|T047|L97.228|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT CALF WITH OTHER SPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF LEFT CALF WITH OTH SEVERITY
C2888674|T047|L97.229|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT CALF WITH UNSPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF LEFT CALF WITH UNSP SEVERITY
C2891204|T037|T85.691A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTRAPERITONEAL DIALYSIS CATHETER, INITIAL ENCOUNTER|MECH COMPL OF INTRAPERITONEAL DIALYSIS CATHETER, INIT ENCNTR
C2888671|T047|L97.222|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT CALF WITH FAT LAYER EXPOSED|NON-PRESSURE CHRONIC ULCER OF LEFT CALF W FAT LAYER EXPOSED
C2888672|T047|L97.223|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT CALF WITH NECROSIS OF MUSCLE|NON-PRESSURE CHRONIC ULCER OF LEFT CALF W NECROSIS OF MUSCLE
C2888670|T047|L97.221|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT CALF LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHRONIC ULCER OF LEFT CALF LIMITED TO BRKDWN SKIN
C4509291|T047|L97.226|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT CALF WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OF LEFT CALF WITH BONE INVL W/O EVD OF NECR
C2888673|T047|L97.224|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT CALF WITH NECROSIS OF BONE|NON-PRESSURE CHRONIC ULCER OF LEFT CALF W NECROSIS OF BONE
C4509290|T047|L97.225|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT CALF WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULCER OF LEFT CALF WITH MSL INVL W/O EVD OF NECR
C0026848|T047|G72.9|DMDICD10|MYOPATHY, UNSPECIFIED|MYOPATHIE, NICHT NAEHER BEZEICHNET
C0410220|T046|G72.0|DMDICD10|DRUG-INDUCED MYOPATHY|ARZNEIMITTELINDUZIERTE MYOPATHIE
C0270985|T047|G72.1|DMDICD10|ALCOHOLIC MYOPATHY|ALKOHOLMYOPATHIE
C0494504|T047|G72.2|DMDICD10|MYOPATHY DUE TO OTHER TOXIC AGENTS|MYOPATHIE DURCH SONSTIGE TOXISCHE AGENZIEN
C2875319|T047|G72.3|ICD10CM|PERIODIC PARALYSIS|NORMOKALEMIC PARALYSIS (FAMILIAL)
C2865561|T037|S88.122S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, LEFT LOWER LEG, SEQUELA|PART TRAUM AMP AT LEVEL BETW KNEE AND ANKLE, L LOW LEG, SQLA
C0263369|T047|L94.5|DMDICD10|POIKILODERMA VASCULARE ATROPHICANS|POIKILODERMIA ATROPHICANS VASCULARIS [JACOBI]
C2874305|T046|E83.32|ICD10CM|HEREDITARY VITAMIN D-DEPENDENT RICKETS (TYPE 1) (TYPE 2)|HEREDITARY VITAMIN D-DEPENDENT RICKETS (TYPE 1) (TYPE 2)
C0494290|T047|E11.9|DMDICD10|TYPE 2 DIABETES MELLITUS WITHOUT COMPLICATIONS|NICHT PRIMAER INSULINABHAENGIGER DIABETES MELLITUS [TYP-II-DIABETES]: OHNE KOMPLIKATIONEN
C1299614|T047|E11.8|DMDICD10|TYPE 2 DIABETES MELLITUS WITH UNSPECIFIED COMPLICATIONS|NICHT PRIMAER INSULINABHAENGIGER DIABETES MELLITUS [TYP-II-DIABETES]: MIT NICHT NAEHER BEZEICHNETEN KOMPLIKATIONEN
C2889049|T047|M02.31|ICD10CM|REITER'S DISEASE, UNSPECIFIED SHOULDER|REITER'S DISEASE, SHOULDER
C2858133|T037|S72.361C|ICD10CM|DISPLACED SEGMENTAL FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL SEG FX SHAFT OF R FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2858132|T037|S72.361B|ICD10CM|DISPLACED SEGMENTAL FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL SEG FX SHAFT OF R FEMUR, INIT FOR OPN FX TYPE I/2
C2858131|T037|S72.361A|ICD10CM|DISPLACED SEGMENTAL FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED SEGMENTAL FRACTURE OF SHAFT OF RIGHT FEMUR, INIT
C2882979|T047|I70.711|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, RIGHT LEG|ATHSCL TYPE OF BYPASS OF THE EXTRM W INTRMT CLAUD, RIGHT LEG
C2889051|T047|M02.312|ICD10CM|REITER'S DISEASE, LEFT SHOULDER|REITER'S DISEASE, LEFT SHOULDER
C2889050|T047|M02.311|ICD10CM|REITER'S DISEASE, RIGHT SHOULDER|REITER'S DISEASE, RIGHT SHOULDER
C2833874|T037|S14.108A|ICD10CM|UNSPECIFIED INJURY AT C8 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY AT C8 LEVEL OF CERVICAL SPINAL CORD, INIT ENCNTR
C0260690|T033|Z93.8|DMDICD10|OTHER ARTIFICIAL OPENING STATUS|VORHANDENSEIN VON SONSTIGEN KUENSTLICHEN KOERPEROEFFNUNGEN
C2876996|T037|T38.0X2A|ICD10CM|POISONING BY GLUCOCORTICOIDS AND SYNTHETIC ANALOGUES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY GLUCOCORT/SYNTH ANALOG, SELF-HARM, INIT
C4290096|T047|E15|ICD10CM|NONDIABETIC HYPOGLYCEMIC COMA|HYPERINSULINISM WITH HYPOGLYCEMIC COMA
C2901816|T047|M86.171|ICD10CM|OTHER ACUTE OSTEOMYELITIS, RIGHT ANKLE AND FOOT|OTHER ACUTE OSTEOMYELITIS, RIGHT ANKLE AND FOOT
C2712692|T191|C4A.4|ICD10CM|MERKEL CELL CARCINOMA OF SCALP AND NECK|MERKEL CELL CARCINOMA OF SCALP AND NECK
C2876998|T037|T38.0X2S|ICD10CM|POISONING BY GLUCOCORTICOIDS AND SYNTHETIC ANALOGUES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY GLUCOCORT/SYNTH ANALOG, SELF-HARM, SEQUELA
C2887058|T047|A31.2|ICD10CM|DISSEMINATED MYCOBACTERIUM AVIUM-INTRACELLULARE COMPLEX (DMAC)|DISSEM MYCOBACTERIUM AVIUM-INTRACELLULARE COMPLEX (DMAC)
C2712673|T191|C4A.0|ICD10CM|MERKEL CELL CARCINOMA OF LIP|MERKEL CELL CARCINOMA OF LIP
C3249882|T047|A31.0|ICD10CM|PULMONARY MYCOBACTERIAL INFECTION|INFECTION DUE TO MYCOBACTERIUM AVIUM
C2837452|T037|S32.001A|ICD10CM|STABLE BURST FRACTURE OF UNSPECIFIED LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|STABLE BURST FRACTURE OF UNSP LUMBAR VERTEBRA, INIT
C2837453|T037|S32.001B|ICD10CM|STABLE BURST FRACTURE OF UNSPECIFIED LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|STABLE BURST FRACTURE OF UNSP LUM VERTEBRA, INIT FOR OPN FX
C2874306|T046|E83.39|ICD10CM|OTHER DISORDERS OF PHOSPHORUS METABOLISM|OTHER DISORDERS OF PHOSPHORUS METABOLISM
C2842074|T191|C4A.8|ICD10CM|MERKEL CELL CARCINOMA OF OVERLAPPING SITES|MERKEL CELL CARCINOMA OF OVERLAPPING SITES
C2977927|T191|C4A.9|ICD10CM|MERKEL CELL CARCINOMA, UNSPECIFIED|MERKEL CELL CARCINOMA OF UNSPECIFIED SITE
C0339009|T048|F91.0|DMDICD10|CONDUCT DISORDER CONFINED TO FAMILY CONTEXT|AUF DEN FAMILIAEREN RAHMEN BESCHRAENKTE STOERUNG DES SOZIALVERHALTENS
C0865417|T048||ICD10CM|CONDUCT DISORDER, CHILDHOOD-ONSET TYPE
C0375192|T048|F91.2|ICD10CM|CONDUCT DISORDER, ADOLESCENT-ONSET TYPE|CONDUCT DISORDER, ADOLESCENT-ONSET TYPE
C0029121|T048|F91.3|DMDICD10|OPPOSITIONAL DEFIANT DISORDER|STOERUNG DES SOZIALVERHALTENS MIT OPPOSITIONELLEM, AUFSAESSIGEM VERHALTEN
C4268307|T048|F91.8|ICD10CM|OTHER CONDUCT DISORDERS|OTHER SPECIFIED DISRUPTIVE DISORDER
C4268308|T048|F91.9|ICD10CM|CONDUCT DISORDER, UNSPECIFIED|DISRUPTIVE DISORDER NOS
C2901818|T047|M86.179|ICD10CM|OTHER ACUTE OSTEOMYELITIS, UNSPECIFIED ANKLE AND FOOT|OTHER ACUTE OSTEOMYELITIS, UNSPECIFIED ANKLE AND FOOT
C2878588|T037|T43.612S|ICD10CM|POISONING BY CAFFEINE, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY CAFFEINE, INTENTIONAL SELF-HARM, SEQUELA
C2853930|T191|C83.58|ICD10CM|LYMPHOBLASTIC (DIFFUSE) LYMPHOMA, LYMPH NODES OF MULTIPLE SITES|LYMPHOBLASTIC (DIFFUSE) LYMPHOMA, LYMPH NODES MULT SITE
C2853931|T191|C83.59|ICD10CM|LYMPHOBLASTIC (DIFFUSE) LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES|LYMPHOBLASTIC LYMPHOMA, EXTRNOD AND SOLID ORGAN SITES
C2893639|T047|M12.039|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], UNSPECIFIED WRIST|CHRONIC POSTRHEUMATIC ARTHROPATHY, UNSPECIFIED WRIST
C2853924|T191|C83.52|ICD10CM|LYMPHOBLASTIC (DIFFUSE) LYMPHOMA, INTRATHORACIC LYMPH NODES|LYMPHOBLASTIC (DIFFUSE) LYMPHOMA, INTRATHORACIC LYMPH NODES
C2853925|T191|C83.53|ICD10CM|LYMPHOBLASTIC (DIFFUSE) LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES|LYMPHOBLASTIC (DIFFUSE) LYMPHOMA, INTRA-ABD LYMPH NODES
C2853922|T191|C83.50|ICD10CM|LYMPHOBLASTIC (DIFFUSE) LYMPHOMA, UNSPECIFIED SITE|LYMPHOBLASTIC (DIFFUSE) LYMPHOMA, UNSPECIFIED SITE
C2853923|T191|C83.51|ICD10CM|LYMPHOBLASTIC (DIFFUSE) LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK|LYMPHOBLASTIC LYMPHOMA, NODES OF HEAD, FACE, AND NECK
C2853928|T191|C83.56|ICD10CM|LYMPHOBLASTIC (DIFFUSE) LYMPHOMA, INTRAPELVIC LYMPH NODES|LYMPHOBLASTIC (DIFFUSE) LYMPHOMA, INTRAPELVIC LYMPH NODES
C2853929|T191|C83.57|ICD10CM|LYMPHOBLASTIC (DIFFUSE) LYMPHOMA, SPLEEN|LYMPHOBLASTIC (DIFFUSE) LYMPHOMA, SPLEEN
C2853926|T191|C83.54|ICD10CM|LYMPHOBLASTIC (DIFFUSE) LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB|LYMPHOBLASTIC LYMPHOMA, NODES OF AXILLA AND UPPER LIMB
C2853927|T191|C83.55|ICD10CM|LYMPHOBLASTIC (DIFFUSE) LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|LYMPHOBLASTIC LYMPHOMA, NODES OF ING REGION AND LOWER LIMB
C2861642|T191|C94.6|ICD10CM|MYELODYSPLASTIC DISEASE, NOT CLASSIFIED|MYELODYSPLASTIC DISEASE, NOT CLASSIFIED
C2877687|T037|T40.5X2A|ICD10CM|POISONING BY COCAINE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY COCAINE, INTENTIONAL SELF-HARM, INIT ENCNTR
C4270469|T046|T85.113A|ICD10CM|BREAKDOWN (MECHANICAL) OF IMPLANTED ELECTRONIC NEUROSTIMULATOR, GENERATOR, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF IMPLNT ELEC NSTIM, GENERATOR, INIT
C2848423|T037|S58.119A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN ELBOW AND WRIST, UNSPECIFIED ARM, INITIAL ENCOUNTER|COMPLETE TRAUM AMP AT LEV BETW ELBOW AND WRS, UNSP ARM, INIT
C2877689|T037|T40.5X2S|ICD10CM|POISONING BY COCAINE, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY COCAINE, INTENTIONAL SELF-HARM, SEQUELA
C2848425|T037|S58.119S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN ELBOW AND WRIST, UNSPECIFIED ARM, SEQUELA|COMPLETE TRAUM AMP AT LEV BETW ELBOW AND WRS, UNSP ARM, SQLA
C2858595|T037|S72.434C|ICD10CM|NONDISPLACED FRACTURE OF MEDIAL CONDYLE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF MED CONDYLE OF R FEMR, 7THC
C0238124|T047|M72.6|ICD10CM|NECROTIZING FASCIITIS|NECROTIZING FASCIITIS
C1571983|T048||ICD10CM|DELUSIONAL DISORDERS
C2888567|T047|L89.621|ICD10CM|PRESSURE ULCER OF LEFT HEEL, STAGE 1|PRESSURE ULCER OF LEFT HEEL, STAGE 1
C2888564|T047||ICD10CM|PRESSURE ULCER OF LEFT HEEL, UNSTAGEABLE
C2888573|T047|L89.623|ICD10CM|PRESSURE ULCER OF LEFT HEEL, STAGE 3|PRESSURE ULCER OF LEFT HEEL, STAGE 3
C2888570|T047|L89.622|ICD10CM|PRESSURE ULCER OF LEFT HEEL, STAGE 2|PRESSURE ULCER OF LEFT HEEL, STAGE 2
C2837589|T037|S32.040A|ICD10CM|WEDGE COMPRESSION FRACTURE OF FOURTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|WEDGE COMPRESSION FRACTURE OF FOURTH LUMBAR VERTEBRA, INIT
C2888579|T047|L89.629|ICD10CM|PRESSURE ULCER OF LEFT HEEL, UNSPECIFIED STAGE|PRESSURE ULCER OF LEFT HEEL, UNSPECIFIED STAGE
C0338590|T047|A52.04|ICD10CM|SYPHILITIC CEREBRAL ARTERITIS|SYPHILITIC CEREBRAL ARTERITIS
C2838634|T037|S34.105S|ICD10CM|UNSPECIFIED INJURY TO L5 LEVEL OF LUMBAR SPINAL CORD, SEQUELA|UNSP INJURY TO L5 LEVEL OF LUMBAR SPINAL CORD, SEQUELA
C2883067|T047|I80.219|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF UNSPECIFIED ILIAC VEIN|PHLEBITIS AND THROMBOPHLEBITIS OF UNSPECIFIED ILIAC VEIN
C2855966|T037|S68.422S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT HAND AT WRIST LEVEL, SEQUELA|PARTIAL TRAUMATIC AMP OF LEFT HAND AT WRIST LEVEL, SEQUELA
C2883064|T047|I80.211|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF RIGHT ILIAC VEIN|PHLEBITIS AND THROMBOPHLEBITIS OF RIGHT ILIAC VEIN
C2883065|T047|I80.212|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF LEFT ILIAC VEIN|PHLEBITIS AND THROMBOPHLEBITIS OF LEFT ILIAC VEIN
C2883066|T047|I80.213|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF ILIAC VEIN, BILATERAL|PHLEBITIS AND THROMBOPHLEBITIS OF ILIAC VEIN, BILATERAL
C2830466|T184|R65.11|ICD10CM|SYSTEMIC INFLAMMATORY RESPONSE SYNDROME (SIRS) OF NON-INFECTIOUS ORIGIN WITH ACUTE ORGAN DYSFUNCTION|SIRS OF NON-INFECTIOUS ORIGIN W ACUTE ORGAN DYSFUNCTION
C2830465|T184|R65.10|ICD10CM|SYSTEMIC INFLAMMATORY RESPONSE SYNDROME (SIRS) OF NON-INFECTIOUS ORIGIN WITHOUT ACUTE ORGAN DYSFUNCTION|SIRS OF NON-INFECTIOUS ORIGIN W/O ACUTE ORGAN DYSFUNCTION
C0153869|T191||ICD10AM|MULTIPLE MYELOMA IN REMISSION
C2854076|T191||ICD10CM|MULTIPLE MYELOMA NOT HAVING ACHIEVED REMISSION
C2887360|T047|I97.810|ICD10CM|INTRAOPERATIVE CEREBROVASCULAR INFARCTION DURING CARDIAC SURGERY|INTRAOPERATIVE CEREBVASC INFARCTION DURING CARDIAC SURGERY
C2349261|T191||ICD10CM|MULTIPLE MYELOMA IN RELAPSE
C2869794|T037|S98.121A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT GREAT TOE, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF RIGHT GREAT TOE, INIT ENCNTR
C2869795|T037|S98.121D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT GREAT TOE, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF RIGHT GREAT TOE, SUBS ENCNTR
C2876235|T037|T32.99|ICD10CM|CORROSIONS INVOLVING 90% OR MORE OF BODY SURFACE WITH 90% OR MORE THIRD DEGREE CORROSION|CORROS 90%/MORE OF BODY SURFC W 90%/MORE THIRD DEGREE CORROS
C0348807|T047|J41.8|DMDICD10|MIXED SIMPLE AND MUCOPURULENT CHRONIC BRONCHITIS|MISCHFORMEN VON EINFACHER UND SCHLEIMIG-EITRIGER CHRONISCHER BRONCHITIS
C0155873|T047|J41.1|DMDICD10|MUCOPURULENT CHRONIC BRONCHITIS|SCHLEIMIG-EITRIGE CHRONISCHE BRONCHITIS
C0155872|T047|J41.0|DMDICD10|SIMPLE CHRONIC BRONCHITIS|EINFACHE CHRONISCHE BRONCHITIS
C2869796|T037|S98.121S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT GREAT TOE, SEQUELA|PARTIAL TRAUMATIC AMPUTATION OF RIGHT GREAT TOE, SEQUELA
C2876228|T037|T32.92|ICD10CM|CORROSIONS INVOLVING 90% OR MORE OF BODY SURFACE WITH 20-29% THIRD DEGREE CORROSION|CORROS 90%/MORE OF BODY SURFACE W 20-29% THIRD DEGREE CORROS
C2876231|T037|T32.95|ICD10CM|CORROSIONS INVOLVING 90% OR MORE OF BODY SURFACE WITH 50-59% THIRD DEGREE CORROSION|CORROS 90%/MORE OF BODY SURFACE W 50-59% THIRD DEGREE CORROS
C2876230|T037|T32.94|ICD10CM|CORROSIONS INVOLVING 90% OR MORE OF BODY SURFACE WITH 40-49% THIRD DEGREE CORROSION|CORROS 90%/MORE OF BODY SURFACE W 40-49% THIRD DEGREE CORROS
C2876233|T037|T32.97|ICD10CM|CORROSIONS INVOLVING 90% OR MORE OF BODY SURFACE WITH 70-79% THIRD DEGREE CORROSION|CORROS 90%/MORE OF BODY SURFACE W 70-79% THIRD DEGREE CORROS
C4236942|T048|F10.96|ICD10CM|ALCOHOL USE, UNSPECIFIED WITH ALCOHOL-INDUCED PERSISTING AMNESTIC DISORDER|ALCOHOL-INDUCED MAJOR NEUROCOGNITIVE DISORDER, AMNESTIC-CONFABULATORY TYPE, WITHOUT USE DISORDER
C2833555|T037|S12.550B|ICD10CM|OTHER TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH TRAUM DISPL SPONDYLOLYSIS OF SIXTH CERVCAL VERT, 7THB
C2833554|T037|S12.550A|ICD10CM|OTHER TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH TRAUM DISPL SPONDYLOLYSIS OF SIXTH CERVCAL VERT, INIT
C2859027|T037|S72.8X1A|ICD10CM|OTHER FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF RIGHT FEMUR, INIT ENCNTR FOR CLOSED FRACTURE
C2859028|T037|S72.8X1B|ICD10CM|OTHER FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|OTH FRACTURE OF RIGHT FEMUR, INIT FOR OPN FX TYPE I/2
C2859029|T037|S72.8X1C|ICD10CM|OTHER FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|OTH FRACTURE OF RIGHT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C0153894|T191|C92.Z1|ICD10CM|OTHER MYELOID LEUKEMIA, IN REMISSION|OTHER MYELOID LEUKEMIA, IN REMISSION
C2861613|T191|C92.Z0|ICD10CM|OTHER MYELOID LEUKEMIA NOT HAVING ACHIEVED REMISSION|OTHER MYELOID LEUKEMIA NOT HAVING ACHIEVED REMISSION
C2833978|T037|S14.136S|ICD10CM|ANTERIOR CORD SYNDROME AT C6 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|ANTERIOR CORD SYNDROME AT C6, SEQUELA
C2349283|T191|C92.Z2|ICD10CM|OTHER MYELOID LEUKEMIA, IN RELAPSE|OTHER MYELOID LEUKEMIA, IN RELAPSE
C2874079|T047|E11.29|ICD10CM|TYPE 2 DIABETES MELLITUS WITH OTHER DIABETIC KIDNEY COMPLICATION|TYPE 2 DIABETES MELLITUS W OTH DIABETIC KIDNEY COMPLICATION
C2876131|T037|T31.21|ICD10CM|BURNS INVOLVING 20-29% OF BODY SURFACE WITH 10-19% THIRD DEGREE BURNS|BURNS OF 20-29% OF BODY SURFACE W 10-19% THIRD DEGREE BURNS
C2874075|T047|E11.21|ICD10CM|TYPE 2 DIABETES MELLITUS WITH DIABETIC NEPHROPATHY|TYPE 2 DIABETES MELLITUS WITH INTRACAPILLARY GLOMERULONEPHROSIS
C2874077|T047|E11.22|ICD10CM|TYPE 2 DIABETES MELLITUS WITH DIABETIC CHRONIC KIDNEY DISEASE|TYPE 2 DIABETES MELLITUS W DIABETIC CHRONIC KIDNEY DISEASE
C2833976|T037|S14.136A|ICD10CM|ANTERIOR CORD SYNDROME AT C6 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|ANTERIOR CORD SYNDROME AT C6, INIT
C2833368|T037|S12.290A|ICD10CM|OTHER DISPLACED FRACTURE OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH DISP FX OF THIRD CERVICAL VERTEBRA, INIT FOR CLOS FX
C2901773|T047|M86.021|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, RIGHT HUMERUS|ACUTE HEMATOGENOUS OSTEOMYELITIS, RIGHT HUMERUS
C2833977|T037|S14.136D|ICD10CM|ANTERIOR CORD SYNDROME AT C6 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|ANTERIOR CORD SYNDROME AT C6, SUBS
C2901774|T047|M86.022|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, LEFT HUMERUS|ACUTE HEMATOGENOUS OSTEOMYELITIS, LEFT HUMERUS
C2901775|T047|M86.029|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED HUMERUS|ACUTE HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED HUMERUS
C2349323|T191||ICD10CM|MALIGNANT CARCINOID TUMOR OF THE SIGMOID COLON
C2349322|T191||ICD10CM|MALIGNANT CARCINOID TUMOR OF THE DESCENDING COLON
C0496944|T191|D44.3|DMDICD10|NEOPLASM OF UNCERTAIN BEHAVIOR OF PITUITARY GLAND|NEUBILDUNG UNSICHEREN ODER UNBEKANNTEN VERHALTENS: HYPOPHYSE
C0496945|T191|D44.4|DMDICD10|NEOPLASM OF UNCERTAIN BEHAVIOR OF CRANIOPHARYNGEAL DUCT|NEUBILDUNG UNSICHEREN ODER UNBEKANNTEN VERHALTENS: DUCTUS CRANIOPHARYNGEALIS
C0496946|T191|D44.5|DMDICD10|NEOPLASM OF UNCERTAIN BEHAVIOR OF PINEAL GLAND|NEUBILDUNG UNSICHEREN ODER UNBEKANNTEN VERHALTENS: EPIPHYSE [GLANDULA PINEALIS] [ZIRBELDRUESE]
C2349321|T191||ICD10CM|MALIGNANT CARCINOID TUMOR OF THE TRANSVERSE COLON
C2349320|T191||ICD10CM|MALIGNANT CARCINOID TUMOR OF THE ASCENDING COLON
C2349318|T191||ICD10CM|MALIGNANT CARCINOID TUMOR OF THE LARGE INTESTINE, UNSPECIFIED PORTION
C2856776|T037|S72.036B|ICD10CM|NONDISPLACED MIDCERVICAL FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP MIDCERVICAL FX UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2856777|T037|S72.036C|ICD10CM|NONDISPLACED MIDCERVICAL FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP MIDCERVICAL FX UNSP FEMR, 7THC
C2856775|T037|S72.036A|ICD10CM|NONDISPLACED MIDCERVICAL FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED MIDCERVICAL FRACTURE OF UNSP FEMUR, INIT
C2842107|T191|C50.419|ICD10CM|MALIGNANT NEOPLASM OF UPPER-OUTER QUADRANT OF UNSPECIFIED FEMALE BREAST|MALIG NEOPLASM OF UPPER-OUTER QUADRANT OF UNSP FEMALE BREAST
C2842105|T191|C50.411|ICD10CM|MALIGNANT NEOPLASM OF UPPER-OUTER QUADRANT OF RIGHT FEMALE BREAST|MALIG NEOPLM OF UPPER-OUTER QUADRANT OF RIGHT FEMALE BREAST
C2842106|T191|C50.412|ICD10CM|MALIGNANT NEOPLASM OF UPPER-OUTER QUADRANT OF LEFT FEMALE BREAST|MALIG NEOPLASM OF UPPER-OUTER QUADRANT OF LEFT FEMALE BREAST
C4269559|T037|S02.672A|ICD10CM|FRACTURE OF ALVEOLUS OF LEFT MANDIBLE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF ALVEOLUS OF LEFT MANDIBLE, INIT
C4269560|T037|S02.672B|ICD10CM|FRACTURE OF ALVEOLUS OF LEFT MANDIBLE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF ALVEOLUS OF LEFT MANDIBLE, 7THB
C2884168|T037|T52.8X2A|ICD10CM|TOXIC EFFECT OF OTHER ORGANIC SOLVENTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF ORGANIC SOLVENTS, SELF-HARM, INIT
C2876770|T037|T36.92XS|ICD10CM|POISONING BY UNSPECIFIED SYSTEMIC ANTIBIOTIC, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY UNSP SYSTEMIC ANTIBIOTIC, SELF-HARM, SEQUELA
C2890068|T037|T82.531A|ICD10CM|LEAKAGE OF SURGICALLY CREATED ARTERIOVENOUS SHUNT, INITIAL ENCOUNTER|LEAKAGE OF SURGICALLY CREATED ARTERIOVENOUS SHUNT, INIT
C2832606|T037|S06.824A|ICD10CM|INJURY OF LEFT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|INJURY OF L INT CAROTID, INTCR W LOC OF 6-24 HRS, INIT
C2888703|T047|L97.411|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT HEEL AND MIDFOOT LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHR ULCER OF RIGHT HEEL AND MIDFT LMT TO BRKDWN SKIN
C2888705|T047|L97.413|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT HEEL AND MIDFOOT WITH NECROSIS OF MUSCLE|NON-PRS CHR ULCER OF RIGHT HEEL AND MIDFOOT W NECROS MUSCLE
C2888704|T047|L97.412|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT HEEL AND MIDFOOT WITH FAT LAYER EXPOSED|NON-PRS CHR ULCER OF RIGHT HEEL AND MIDFT W FAT LAYER EXPOS
C4509305|T047|L97.415|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT HEEL AND MIDFOOT WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OF R HEEL/MIDFT W MSL INVL W/O EVD OF NECR
C2888706|T047|L97.414|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT HEEL AND MIDFOOT WITH NECROSIS OF BONE|NON-PRS CHR ULCER OF RIGHT HEEL AND MIDFOOT W NECROS BONE
C4509306|T047|L97.416|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT HEEL AND MIDFOOT WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OF R HEEL/MIDFT W BNE INVL W/O EVD OF NECR
C2888707|T047|L97.419|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT HEEL AND MIDFOOT WITH UNSPECIFIED SEVERITY|NON-PRS CHR ULCER OF RIGHT HEEL AND MIDFOOT W UNSP SEVERT
C2889012|T047|M02.159|ICD10CM|POSTDYSENTERIC ARTHROPATHY, UNSPECIFIED HIP|POSTDYSENTERIC ARTHROPATHY, UNSPECIFIED HIP
C2895358|T047|M49.87|ICD10CM|SPONDYLOPATHY IN DISEASES CLASSIFIED ELSEWHERE, LUMBOSACRAL REGION|SPONDYLOPATHY IN DISEASES CLASSD ELSWHR, LUMBOSACRAL REGION
C2895357|T047|M49.86|ICD10CM|SPONDYLOPATHY IN DISEASES CLASSIFIED ELSEWHERE, LUMBAR REGION|SPONDYLOPATHY IN DISEASES CLASSD ELSWHR, LUMBAR REGION
C2895352|T047|M49.81|ICD10CM|SPONDYLOPATHY IN DISEASES CLASSIFIED ELSEWHERE, OCCIPITO-ATLANTO-AXIAL REGION|SPOND IN DISEASES CLASSD ELSWHR, OCCIPT-ATLAN-AX REGION
C2895351|T047|M49.80|ICD10CM|SPONDYLOPATHY IN DISEASES CLASSIFIED ELSEWHERE, SITE UNSPECIFIED|SPONDYLOPATHY IN DISEASES CLASSIFIED ELSEWHERE, SITE UNSP
C2895354|T047|M49.83|ICD10CM|SPONDYLOPATHY IN DISEASES CLASSIFIED ELSEWHERE, CERVICOTHORACIC REGION|SPONDYLOPATHY IN DISEASES CLASSD ELSWHR, CERVICOTHOR REGION
C2895353|T047|M49.82|ICD10CM|SPONDYLOPATHY IN DISEASES CLASSIFIED ELSEWHERE, CERVICAL REGION|SPONDYLOPATHY IN DISEASES CLASSD ELSWHR, CERVICAL REGION
C2883120|T047|I82.511|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF RIGHT FEMORAL VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF RIGHT FEMORAL VEIN
C0839986|T047||ICD10AM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, OTHER SITE
C2883122|T047|I82.513|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF FEMORAL VEIN, BILATERAL|CHRONIC EMBOLISM AND THROMBOSIS OF FEMORAL VEIN, BILATERAL
C2883121|T047|I82.512|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF LEFT FEMORAL VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF LEFT FEMORAL VEIN
C2883123|T047|I82.519|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED FEMORAL VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED FEMORAL VEIN
C0839978|T047||ICD10AM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED SITE
C2890588|T037|T84.112A|ICD10CM|BREAKDOWN (MECHANICAL) OF INTERNAL FIXATION DEVICE OF BONE OF RIGHT FOREARM, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF INT FIX OF BONE OF R FOREARM, INIT
C2889211|T047|M05.339|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP WRIST
C2833852|T037|S14.102S|ICD10CM|UNSPECIFIED INJURY AT C2 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|UNSP INJURY AT C2 LEVEL OF CERVICAL SPINAL CORD, SEQUELA
C2893328|T047|A50.55|ICD10CM|LATE CONGENITAL SYPHILITIC ARTHROPATHY|LATE CONGENITAL SYPHILITIC ARTHROPATHY
C2889210|T047|M05.332|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT WRIST|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF L WRIST
C2879671|T037|T47.0X2A|ICD10CM|POISONING BY HISTAMINE H2-RECEPTOR BLOCKERS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY HISTAMINE H2-RECEPTOR BLOCKERS, SELF-HARM, INIT
C2889079|T047|M02.811|ICD10CM|OTHER REACTIVE ARTHROPATHIES, RIGHT SHOULDER|OTHER REACTIVE ARTHROPATHIES, RIGHT SHOULDER
C2889080|T047|M02.812|ICD10CM|OTHER REACTIVE ARTHROPATHIES, LEFT SHOULDER|OTHER REACTIVE ARTHROPATHIES, LEFT SHOULDER
C2889010|T047|M02.151|ICD10CM|POSTDYSENTERIC ARTHROPATHY, RIGHT HIP|POSTDYSENTERIC ARTHROPATHY, RIGHT HIP
C2937222|T047||ICD10CM|ULCERATIVE (CHRONIC) PROCTITIS WITHOUT COMPLICATIONS
C2889078|T047|M02.81|ICD10CM|OTHER REACTIVE ARTHROPATHIES, UNSPECIFIED SHOULDER|OTHER REACTIVE ARTHROPATHIES, SHOULDER
C2874267|T047|E74.09|ICD10CM|OTHER GLYCOGEN STORAGE DISEASE|OTHER GLYCOGEN STORAGE DISEASE
C2902080|T046|M87.30|ICD10CM|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED BONE|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED BONE
C3264595|T048|F40.02|ICD10CM|AGORAPHOBIA WITHOUT PANIC DISORDER|AGORAPHOBIA WITHOUT PANIC DISORDER
C0236800|T048||ICD10AM|AGORAPHOBIA WITH PANIC DISORDER
C0001819|T048|F40.00|ICD10AM|AGORAPHOBIA, UNSPECIFIED|AGORAPHOBIA WITHOUT MENTION OF PANIC DISORDER
C0017920|T047||ICD10CM|VON GIERKE DISEASE
C0017919|T047|E74.00|ICD10CM|GLYCOGEN STORAGE DISEASE, UNSPECIFIED|GLYCOGEN STORAGE DISEASE, UNSPECIFIED
C0017922|T047||ICD10CM|CORI DISEASE
C0155998|T047|K26.2|DMDICD10|ACUTE DUODENAL ULCER WITH BOTH HEMORRHAGE AND PERFORATION|ULCUS DUODENI: AKUT, MIT BLUTUNG UND PERFORATION
C0391983|T047|K26.5|DMDICD10|CHRONIC OR UNSPECIFIED DUODENAL ULCER WITH PERFORATION|ULCUS DUODENI: CHRONISCH ODER NICHT NAEHER BEZEICHNET, MIT PERFORATION
C0017924|T047||ICD10CM|MCARDLE DISEASE
C0494726|T047|K26.6|DMDICD10|CHRONIC OR UNSPECIFIED DUODENAL ULCER WITH BOTH HEMORRHAGE AND PERFORATION|ULCUS DUODENI: CHRONISCH ODER NICHT NAEHER BEZEICHNET, MIT BLUTUNG UND PERFORATION
C2883889|T037|T50.B12S|ICD10CM|POISONING BY SMALLPOX VACCINES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY SMALLPOX VACCINES, SELF-HARM, SEQUELA
C2838651|T037|S34.113S|ICD10CM|COMPLETE LESION OF L3 LEVEL OF LUMBAR SPINAL CORD, SEQUELA|COMPLETE LESION OF L3 LEVEL OF LUMBAR SPINAL CORD, SEQUELA
C2901117|T046|M84.479A|ICD10CM|PATHOLOGICAL FRACTURE, UNSPECIFIED TOE(S), INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, UNSP TOE(S), INIT ENCNTR FOR FRACTURE
C0694507|T047|K67|DMDICD10|DISORDERS OF PERITONEUM IN INFECTIOUS DISEASES CLASSIFIED ELSEWHERE|KRANKHEITEN DES PERITONEUMS BEI ANDERENORTS KLASSIFIZIERTEN INFEKTIONSKRANKHEITEN
C2838649|T037|S34.113A|ICD10CM|COMPLETE LESION OF L3 LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION OF L3 LEVEL OF LUMBAR SPINAL CORD, INIT
C2838650|T037|S34.113D|ICD10CM|COMPLETE LESION OF L3 LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION OF L3 LEVEL OF LUMBAR SPINAL CORD, SUBS
C2887101|T047|A41.9|ICD10CM|SEPSIS, UNSPECIFIED ORGANISM|SEPSIS, UNSPECIFIED ORGANISM
C2885285|T037|T62.92XA|ICD10CM|TOXIC EFFECT OF UNSPECIFIED NOXIOUS SUBSTANCE EATEN AS FOOD, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFF OF UNSP NOXIOUS SUB EATEN AS FOOD, SLF-HRM, INIT
C2887089|T047|A41.1|ICD10CM|SEPSIS DUE TO OTHER SPECIFIED STAPHYLOCOCCUS|SEPSIS DUE TO OTHER SPECIFIED STAPHYLOCOCCUS
C2887090|T047|A41.2|ICD10CM|SEPSIS DUE TO UNSPECIFIED STAPHYLOCOCCUS|SEPSIS DUE TO UNSPECIFIED STAPHYLOCOCCUS
C2887091|T047||ICD10CM|SEPSIS DUE TO HEMOPHILUS INFLUENZAE
C2887092|T047|A41.4|ICD10CM|SEPSIS DUE TO ANAEROBES|SEPSIS DUE TO ANAEROBES
C2885287|T037|T62.92XS|ICD10CM|TOXIC EFFECT OF UNSPECIFIED NOXIOUS SUBSTANCE EATEN AS FOOD, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFF OF UNSP NOXIOUS SUB EATEN AS FOOD, SLF-HRM, SQLA
C2832180|T037|S06.330S|ICD10CM|CONTUSION AND LACERATION OF CEREBRUM, UNSPECIFIED, WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|CONTUS/LAC CEREB, W/O LOSS OF CONSCIOUSNESS, SEQUELA
C0282528|T047|E71.50|ICD10CM|PEROXISOMAL DISORDER, UNSPECIFIED|PEROXISOMAL DISORDER, UNSPECIFIED
C2875047|T047|G11.3|ICD10CM|CEREBELLAR ATAXIA WITH DEFECTIVE DNA REPAIR|ATAXIA TELANGIECTASIA [LOUIS-BAR]
C0393524|T047|G11.2|DMDICD10|LATE-ONSET CEREBELLAR ATAXIA|SPAET BEGINNENDE ZEREBELLARE ATAXIE
C2875046|T047|G11.1|ICD10CM|EARLY-ONSET CEREBELLAR ATAXIA|X-LINKED RECESSIVE SPINOCEREBELLAR ATAXIA
C0394004|T047|G11.0|DMDICD10|CONGENITAL NONPROGRESSIVE ATAXIA|ANGEBORENE NICHTPROGRESSIVE ATAXIE
C2878509|T037|T43.502A|ICD10CM|POISONING BY UNSPECIFIED ANTIPSYCHOTICS AND NEUROLEPTICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY UNSP ANTIPSYCHOT/NEUROLEPT, SELF-HARM, INIT
C4509262|T047|K56.609|ICD10CM|UNSPECIFIED INTESTINAL OBSTRUCTION, UNSPECIFIED AS TO PARTIAL VERSUS COMPLETE OBSTRUCTION|UNSP INTESTNL OBST, UNSP AS TO PARTIAL VERSUS COMPLETE OBST
C2875049|T047|G11.9|ICD10CM|HEREDITARY ATAXIA, UNSPECIFIED|HEREDITARY CEREBELLAR SYNDROME
C0477348|T047|G11.8|DMDICD10|OTHER HEREDITARY ATAXIAS|SONSTIGE HEREDITAERE ATAXIEN
C4509260|T047|K56.600|ICD10CM|PARTIAL INTESTINAL OBSTRUCTION, UNSPECIFIED AS TO CAUSE|INCOMPLETE INTESTINAL OBSTRUCTION, NOS
C4509261|T047|K56.601|ICD10CM|COMPLETE INTESTINAL OBSTRUCTION, UNSPECIFIED AS TO CAUSE|COMPLETE INTESTINAL OBSTRUCTION, UNSPECIFIED AS TO CAUSE
C2873770|T047|D57.80|ICD10CM|OTHER SICKLE-CELL DISORDERS WITHOUT CRISIS|OTHER SICKLE-CELL DISORDERS WITHOUT CRISIS
C2887415|T047|J15.29|ICD10CM|PNEUMONIA DUE TO OTHER STAPHYLOCOCCUS|PNEUMONIA DUE TO OTHER STAPHYLOCOCCUS
C2878511|T037|T43.502S|ICD10CM|POISONING BY UNSPECIFIED ANTIPSYCHOTICS AND NEUROLEPTICS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY UNSP ANTIPSYCHOT/NEUROLEPT, SELF-HARM, SEQUELA
C0032308|T047|J15.20|ICD10CM|PNEUMONIA DUE TO STAPHYLOCOCCUS, UNSPECIFIED|PNEUMONIA DUE TO STAPHYLOCOCCUS, UNSPECIFIED
C2902146|T046|M87.844|ICD10CM|OTHER OSTEONECROSIS, RIGHT FINGER(S)|OTHER OSTEONECROSIS, RIGHT FINGER(S)
C2902147|T046|M87.845|ICD10CM|OTHER OSTEONECROSIS, LEFT FINGER(S)|OTHER OSTEONECROSIS, LEFT FINGER(S)
C4269459|T037|S02.612S|ICD10CM|FRACTURE OF CONDYLAR PROCESS OF LEFT MANDIBLE, SEQUELA|FRACTURE OF CONDYLAR PROCESS OF LEFT MANDIBLE, SEQUELA
C2902143|T046|M87.841|ICD10CM|OTHER OSTEONECROSIS, RIGHT HAND|OTHER OSTEONECROSIS, RIGHT HAND
C2902144|T046|M87.842|ICD10CM|OTHER OSTEONECROSIS, LEFT HAND|OTHER OSTEONECROSIS, LEFT HAND
C2902145|T046|M87.843|ICD10CM|OTHER OSTEONECROSIS, UNSPECIFIED HAND|OTHER OSTEONECROSIS, UNSPECIFIED HAND
C2885407|T037|T63.072A|ICD10CM|TOXIC EFFECT OF VENOM OF OTHER AUSTRALIAN SNAKE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF AUSTRALIAN SNAKE, SELF-HARM, INIT
C2848436|T037|S58.129A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN ELBOW AND WRIST, UNSPECIFIED ARM, INITIAL ENCOUNTER|PART TRAUM AMP AT LEVEL BETW ELBOW AND WRIST, UNSP ARM, INIT
C2902148|T046|M87.849|ICD10CM|OTHER OSTEONECROSIS, UNSPECIFIED FINGER(S)|OTHER OSTEONECROSIS, UNSPECIFIED FINGER(S)
C2835443|T037|S22.080B|ICD10CM|WEDGE COMPRESSION FRACTURE OF T11-T12 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|WEDGE COMPRSN FRACTURE OF T11-T12 VERTEBRA, INIT FOR OPN FX
C0154706|T047|G83.89|ICD10CM|OTHER SPECIFIED PARALYTIC SYNDROMES|OTHER SPECIFIED PARALYTIC SYNDROMES
C2837860|T037|S32.316A|ICD10CM|NONDISPLACED AVULSION FRACTURE OF UNSPECIFIED ILIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED AVULSION FRACTURE OF UNSP ILIUM, INIT
C2883101|T047|I82.429|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED ILIAC VEIN|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED ILIAC VEIN
C4269455|T037|S02.612B|ICD10CM|FRACTURE OF CONDYLAR PROCESS OF LEFT MANDIBLE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF CONDYLAR PROCESS OF LEFT MANDIBLE, 7THB
C4269454|T037|S02.612A|ICD10CM|FRACTURE OF CONDYLAR PROCESS OF LEFT MANDIBLE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF CONDYLAR PROCESS OF LEFT MANDIBLE, INIT
C0242644|T047||ICD10CM|BROWN-SEQUARD SYNDROME
C1859726|T047||ICD10CM|ARTERIAL TORTUOSITY SYNDROME
C0560650|T037|G83.83|ICD10CM|POSTERIOR CORD SYNDROME|POSTERIOR CORD SYNDROME
C0560649|T037|G83.82|ICD10CM|ANTERIOR CORD SYNDROME|ANTERIOR CORD SYNDROME
C2875358|T047|G83.84|ICD10CM|TODD'S PARALYSIS (POSTEPILEPTIC)|TODD'S PARALYSIS (POSTEPILEPTIC)
C2848438|T037|S58.129S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN ELBOW AND WRIST, UNSPECIFIED ARM, SEQUELA|PART TRAUM AMP AT LEVEL BETW ELBOW AND WRIST, UNSP ARM, SQLA
C2856103|T037|S68.722A|ICD10CM|PARTIAL TRAUMATIC TRANSMETACARPAL AMPUTATION OF LEFT HAND, INITIAL ENCOUNTER|PARTIAL TRAUMATIC TRANSMETCRPL AMPUTATION OF LEFT HAND, INIT
C0155626|T047|I21.9|DMDICD10|ACUTE MYOCARDIAL INFARCTION, UNSPECIFIED|AKUTER MYOKARDINFARKT, NICHT NAEHER BEZEICHNET
C4509199|T047|I21.3|ICD10CM|ST ELEVATION (STEMI) MYOCARDIAL INFARCTION OF UNSPECIFIED SITE|TYPE 1 ST ELEVATION MYOCARDIAL INFARCTION OF UNSPECIFIED SITE
C4509200|T047|I21.4|ICD10CM|NON-ST ELEVATION (NSTEMI) MYOCARDIAL INFARCTION|TYPE 1 NON-ST ELEVATION MYOCARDIAL INFARCTION
C2856105|T037|S68.722S|ICD10CM|PARTIAL TRAUMATIC TRANSMETACARPAL AMPUTATION OF LEFT HAND, SEQUELA|PARTIAL TRAUMATIC TRANSMETCRPL AMP OF LEFT HAND, SEQUELA
C2889490|T047|M06.872|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, LEFT ANKLE AND FOOT|OTHER SPECIFIED RHEUMATOID ARTHRITIS, LEFT ANKLE AND FOOT
C2857651|T037|S72.26XC|ICD10CM|NONDISPLACED SUBTROCHANTERIC FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP SUBTROCHNT FX UNSP FEMR, INIT FOR OPN FX TYPE 3A/B/C
C2857650|T037|S72.26XB|ICD10CM|NONDISPLACED SUBTROCHANTERIC FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP SUBTROCHNT FX UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2857649|T037|S72.26XA|ICD10CM|NONDISPLACED SUBTROCHANTERIC FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED SUBTROCHANTERIC FRACTURE OF UNSP FEMUR, INIT
C2877175|T037|T38.7X2S|ICD10CM|POISONING BY ANDROGENS AND ANABOLIC CONGENERS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY ANDROGENS AND ANABOLIC CONGENERS, SLF-HRM, SEQUELA
C2889489|T047|M06.871|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, RIGHT ANKLE AND FOOT|OTHER SPECIFIED RHEUMATOID ARTHRITIS, RIGHT ANKLE AND FOOT
C2837990|T191|C43.22|ICD10CM|MALIGNANT MELANOMA OF LEFT EAR AND EXTERNAL AURICULAR CANAL|MALIGNANT MELANOMA OF LEFT EAR AND EXTERNAL AURICULAR CANAL
C2837989|T191|C43.21|ICD10CM|MALIGNANT MELANOMA OF RIGHT EAR AND EXTERNAL AURICULAR CANAL|MALIGNANT MELANOMA OF RIGHT EAR AND EXTERNAL AURICULAR CANAL
C2837988|T191|C43.20|ICD10CM|MALIGNANT MELANOMA OF UNSPECIFIED EAR AND EXTERNAL AURICULAR CANAL|MALIGNANT MELANOMA OF UNSP EAR AND EXTERNAL AURICULAR CANAL
C2887283|T047|I87.031|ICD10CM|POSTTHROMBOTIC SYNDROME WITH ULCER AND INFLAMMATION OF RIGHT LOWER EXTREMITY|POSTTHROM SYNDROME W ULCER AND INFLAMMATION OF R LOW EXTREM
C2887285|T047|I87.033|ICD10CM|POSTTHROMBOTIC SYNDROME WITH ULCER AND INFLAMMATION OF BILATERAL LOWER EXTREMITY|POSTTHROM SYNDROME W ULCER AND INFLAM OF BILATERAL LOW EXTRM
C2887284|T047|I87.032|ICD10CM|POSTTHROMBOTIC SYNDROME WITH ULCER AND INFLAMMATION OF LEFT LOWER EXTREMITY|POSTTHROM SYNDROME W ULCER AND INFLAMMATION OF L LOW EXTREM
C4267941|T047|E08.3551|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, RIGHT EYE|DIABETES WITH STABLE PROLIF DIABETIC RETINOPATHY, RIGHT EYE
C4267943|T047|E08.3553|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, BILATERAL|DIABETES WITH STABLE PROLIF DIABETIC RETINOPATHY, BILATERAL
C4267942|T047|E08.3552|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, LEFT EYE|DIABETES WITH STABLE PROLIF DIABETIC RETINOPATHY, LEFT EYE
C2887286|T047|I87.039|ICD10CM|POSTTHROMBOTIC SYNDROME WITH ULCER AND INFLAMMATION OF UNSPECIFIED LOWER EXTREMITY|POSTTHROM SYNDROME W ULCER AND INFLAM OF UNSP LOW EXTRM
C4267944|T047|E08.3559|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, UNSPECIFIED EYE|DIABETES WITH STABLE PROLIF DIABETIC RETINOPATHY, UNSP
C2889390|T047|M06.01|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, UNSPECIFIED SHOULDER|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, SHOULDER
C2843323|T037|S48.911S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT SHOULDER AND UPPER ARM, LEVEL UNSPECIFIED, SEQUELA|COMPLETE TRAUM AMP OF RIGHT SHLDR/UP ARM, LEVEL UNSP, SQLA
C2889388|T047|M06.011|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, RIGHT SHOULDER|RHEUMATOID ARTHRITIS W/O RHEUMATOID FACTOR, RIGHT SHOULDER
C2889389|T047|M06.012|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, LEFT SHOULDER|RHEUMATOID ARTHRITIS W/O RHEUMATOID FACTOR, LEFT SHOULDER
C2878226|T037|T42.72XA|ICD10CM|POISONING BY UNSPECIFIED ANTIEPILEPTIC AND SEDATIVE-HYPNOTIC DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY UNSP ANTIEPLPTC AND SED-HYPNTC DRUGS, SLF-HRM, INIT
C2878228|T037|T42.72XS|ICD10CM|POISONING BY UNSPECIFIED ANTIEPILEPTIC AND SEDATIVE-HYPNOTIC DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY UNSP ANTIEPLPTC AND SED-HYPNTC DRUGS, SLF-HRM, SQLA
C4237081|T048|F14.959|ICD10CM|COCAINE USE, UNSPECIFIED WITH COCAINE-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|COCAINE INDUCED PSYCHOTIC DISORDER, WITHOUT USE DISORDER
C2890914|T037|T84.85XA|ICD10CM|STENOSIS DUE TO INTERNAL ORTHOPEDIC PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|STENOSIS DUE TO INTERNAL ORTHOPEDIC PROSTH DEV/GRFT, INIT
C2856708|T037|S72.032B|ICD10CM|DISPLACED MIDCERVICAL FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPLACED MIDCERVICAL FX L FEMUR, INIT FOR OPN FX TYPE I/2
C2874616|T048|F14.951|ICD10CM|COCAINE USE, UNSPECIFIED WITH COCAINE-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|COCAINE USE, UNSP W COCAINE-INDUC PSYCH DISORDER W HALLUCIN
C2874615|T048|F14.950|ICD10CM|COCAINE USE, UNSPECIFIED WITH COCAINE-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|COCAINE USE, UNSP W COCAINE-INDUC PSYCH DISORDER W DELUSIONS
C2856709|T037|S72.032C|ICD10CM|DISPLACED MIDCERVICAL FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL MIDCERVICAL FX L FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2856707|T037|S72.032A|ICD10CM|DISPLACED MIDCERVICAL FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED MIDCERVICAL FRACTURE OF LEFT FEMUR, INIT
C0153693|T191|C79.82|ICD10AM|SECONDARY MALIGNANT NEOPLASM OF GENITAL ORGANS|SECONDARY MALIGNANT NEOPLASM OF GENITAL ORGANS
C0346993|T191|C79.81|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF BREAST|SECONDARY MALIGNANT NEOPLASM OF BREAST
C2886753|T037|T79.A11A|ICD10CM|TRAUMATIC COMPARTMENT SYNDROME OF RIGHT UPPER EXTREMITY, INITIAL ENCOUNTER|TRAUMATIC COMPARTMENT SYNDROME OF R UP EXTREM, INIT
C0153684|T191|C79.8|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF OTHER SPECIFIED SITES|SECONDARY MALIGNANT NEOPLASM OF OTHER SPECIFIED SITES
C2832264|T037|S06.350S|ICD10CM|TRAUMATIC HEMORRHAGE OF LEFT CEREBRUM WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|TRAUM HEMOR LEFT CEREBRUM W/O LOSS OF CONSCIOUSNESS, SEQUELA
C2890234|T037|T83.090A|ICD10CM|OTHER MECHANICAL COMPLICATION OF CYSTOSTOMY CATHETER, INITIAL ENCOUNTER|MECH COMPL OF CYSTOSTOMY CATHETER, INITIAL ENCOUNTER
C2860104|T037|S79.092A|ICD10CM|OTHER PHYSEAL FRACTURE OF UPPER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH PHYSEAL FRACTURE OF UPPER END OF LEFT FEMUR, INIT
C0030299|T047|K86.3|DMDICD10|PSEUDOCYST OF PANCREAS|PSEUDOZYSTE DES PANKREAS
C0030283|T047|K86.2|DMDICD10|CYST OF PANCREAS|PANKREASZYSTE
C2074913|T047||ICD10CM|OTHER CHRONIC PANCREATITIS
C0341470|T047|K86.0|DMDICD10|ALCOHOL-INDUCED CHRONIC PANCREATITIS|ALKOHOLINDUZIERTE CHRONISCHE PANKREATITIS
C2901826|T047|M86.231|ICD10CM|SUBACUTE OSTEOMYELITIS, RIGHT RADIUS AND ULNA|SUBACUTE OSTEOMYELITIS, RIGHT RADIUS AND ULNA
C0030286|T047|K86.9|DMDICD10|DISEASE OF PANCREAS, UNSPECIFIED|KRANKHEIT DES PANKREAS, NICHT NAEHER BEZEICHNET
C2842099|T191|C50.312|ICD10CM|MALIGNANT NEOPLASM OF LOWER-INNER QUADRANT OF LEFT FEMALE BREAST|MALIG NEOPLASM OF LOWER-INNER QUADRANT OF LEFT FEMALE BREAST
C2842098|T191|C50.311|ICD10CM|MALIGNANT NEOPLASM OF LOWER-INNER QUADRANT OF RIGHT FEMALE BREAST|MALIG NEOPLM OF LOWER-INNER QUADRANT OF RIGHT FEMALE BREAST
C0037926|T047||ICD10CM|UNSPECIFIED CORD COMPRESSION
C2873945|T047|E08.69|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH OTHER SPECIFIED COMPLICATION|DIABETES DUE TO UNDERLYING CONDITION W OTH COMPLICATION
C0154035|T191|D32.1|DMDICD10|BENIGN NEOPLASM OF SPINAL MENINGES|GUTARTIGE NEUBILDUNG: RUECKENMARKHAEUTE
C0154033|T191|D32.0|DMDICD10|BENIGN NEOPLASM OF CEREBRAL MENINGES|GUTARTIGE NEUBILDUNG: HIRNHAEUTE
C2873944|T047|E08.65|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH HYPERGLYCEMIA|DIABETES DUE TO UNDERLYING CONDITION W HYPERGLYCEMIA
C2875389|T047|G95.29|ICD10CM|OTHER CORD COMPRESSION|OTHER CORD COMPRESSION
C0393847|T047|G61.82|ICD10CM|MULTIFOCAL MOTOR NEUROPATHY|MMN
C0477393|T047|G61.8|ICD10CM|OTHER INFLAMMATORY POLYNEUROPATHIES|OTHER INFLAMMATORY POLYNEUROPATHIES
C3263975|T047|G40.802|ICD10CM|OTHER EPILEPSY, NOT INTRACTABLE, WITHOUT STATUS EPILEPTICUS|OTHER EPILEPSY, NOT INTRACTABLE, WITHOUT STATUS EPILEPTICUS
C2902369|T047|M89.641|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, RIGHT HAND|OSTEOPATHY AFTER POLIOMYELITIS, RIGHT HAND
C2902370|T047|M89.642|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, LEFT HAND|OSTEOPATHY AFTER POLIOMYELITIS, LEFT HAND
C4268017|T047|E10.3293|ICD10CM|TYPE 1 DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|TYPE 1 DIAB WITH MILD NONP RTNOP WITHOUT MACULAR EDEMA, BI
C2889638|T047|M08.941|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, RIGHT HAND|JUVENILE ARTHRITIS, UNSPECIFIED, RIGHT HAND
C2889639|T047|M08.942|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, LEFT HAND|JUVENILE ARTHRITIS, UNSPECIFIED, LEFT HAND
C2891327|T037|T87.33|ICD10CM|NEUROMA OF AMPUTATION STUMP, RIGHT LOWER EXTREMITY|NEUROMA OF AMPUTATION STUMP, RIGHT LOWER EXTREMITY
C2891326|T037|T87.32|ICD10CM|NEUROMA OF AMPUTATION STUMP, LEFT UPPER EXTREMITY|NEUROMA OF AMPUTATION STUMP, LEFT UPPER EXTREMITY
C2891325|T037|T87.31|ICD10CM|NEUROMA OF AMPUTATION STUMP, RIGHT UPPER EXTREMITY|NEUROMA OF AMPUTATION STUMP, RIGHT UPPER EXTREMITY
C2886879|T037|T81.502D|ICD10CM|UNSPECIFIED COMPLICATION OF FOREIGN BODY ACCIDENTALLY LEFT IN BODY FOLLOWING KIDNEY DIALYSIS, SUBSEQUENT ENCOUNTER|UNSP COMP OF FB ACC LEFT IN BODY FOL KIDNEY DIALYSIS, SUBS
C2891328|T037|T87.34|ICD10CM|NEUROMA OF AMPUTATION STUMP, LEFT LOWER EXTREMITY|NEUROMA OF AMPUTATION STUMP, LEFT LOWER EXTREMITY
C0002881|T019|D58.9|DMDICD10|HEREDITARY HEMOLYTIC ANEMIA, UNSPECIFIED|HEREDITAERE HAEMOLYTISCHE ANAEMIE, NICHT NAEHER BEZEICHNET
C0272048|T047|D58.8|ICD10CM|OTHER SPECIFIED HEREDITARY HEMOLYTIC ANEMIAS|STOMATOCYTOSIS
C2884020|T037|T51.2X2S|ICD10CM|TOXIC EFFECT OF 2-PROPANOL, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF 2-PROPANOL, INTENTIONAL SELF-HARM, SEQUELA
C2831988|T037|S06.1X4A|ICD10CM|TRAUMATIC CEREBRAL EDEMA WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|TRAUMATIC CEREBRAL EDEMA W LOC OF 6 HOURS TO 24 HOURS, INIT
C4268018|T047|E10.3299|ICD10CM|TYPE 1 DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|TYPE 1 DIAB WITH MILD NONP RTNOP WITHOUT MACULAR EDEMA, UNSP
C0013902|T047|D58.1|DMDICD10|HEREDITARY ELLIPTOCYTOSIS|HEREDITAERE ELLIPTOZYTOSE
C2873774|T047|D58.0|ICD10CM|HEREDITARY SPHEROCYTOSIS|CONGENITAL (SPHEROCYTIC) HEMOLYTIC ICTERUS
C0272080|T047||ICD10CM|OTHER HEMOGLOBINOPATHIES
C0494514|T046|G93.1|DMDICD10|ANOXIC BRAIN DAMAGE, NOT ELSEWHERE CLASSIFIED|ANOXISCHE HIRNSCHAEDIGUNG, ANDERENORTS NICHT KLASSIFIZIERT
C2910848|T033|Z44.129|ICD10CM|ENCOUNTER FOR FITTING AND ADJUSTMENT OF PARTIAL ARTIFICIAL LEG, UNSPECIFIED LEG|ENCOUNTER FOR FIT/ADJST OF PARTIAL ARTIFICIAL LEG, UNSP LEG
C2875381|T047|G93.5|ICD10CM|COMPRESSION OF BRAIN|ARNOLD-CHIARI TYPE 1 COMPRESSION OF BRAIN
C2874495|T048|F12.29|ICD10CM|CANNABIS DEPENDENCE WITH UNSPECIFIED CANNABIS-INDUCED DISORDER|CANNABIS DEPENDENCE WITH UNSP CANNABIS-INDUCED DISORDER
C0035400|T047|G93.7|DMDICD10|REYE'S SYNDROME|REYE-SYNDROM
C0006114|T047|G93.6|DMDICD10|CEREBRAL EDEMA|HIRNOEDEM
C2910847|T033|Z44.122|ICD10CM|ENCOUNTER FOR FITTING AND ADJUSTMENT OF PARTIAL ARTIFICIAL LEFT LEG|ENCOUNTER FOR FIT/ADJST OF PARTIAL ARTIFICIAL LEFT LEG
C2831990|T037|S06.1X4S|ICD10CM|TRAUMATIC CEREBRAL EDEMA WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|TRAUMATIC CEREBRAL EDEMA W LOC OF 6-24 HRS, SEQUELA
C4237028|T048|F12.20|ICD10CM|CANNABIS DEPENDENCE, UNCOMPLICATED|CANNABIS USE DISORDER, SEVERE
C4509049|T048|F12.21|ICD10CM|CANNABIS DEPENDENCE, IN REMISSION|CANNABIS USE DISORDER, SEVERE, IN SUSTAINED REMISSION
C2874007|T047|E09.630|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PERIODONTAL DISEASE|DRUG/CHEM DIABETES MELLITUS W PERIODONTAL DISEASE
C2905673|T037|X72.XXXD|ICD10CM|INTENTIONAL SELF-HARM BY HANDGUN DISCHARGE, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY HANDGUN DISCHARGE, SUBS ENCNTR
C4269336|T037|S02.30XB|ICD10CM|FRACTURE OF ORBITAL FLOOR, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF ORBITAL FLOOR, UNSPECIFIED SIDE, 7THB
C4269335|T037|S02.30XA|ICD10CM|FRACTURE OF ORBITAL FLOOR, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF ORBITAL FLOOR, UNSPECIFIED SIDE, INIT
C2877739|T037|T40.692A|ICD10CM|POISONING BY OTHER NARCOTICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH NARCOTICS, INTENTIONAL SELF-HARM, INIT
C2859194|T037|S73.023A|ICD10CM|OBTURATOR SUBLUXATION OF UNSPECIFIED HIP, INITIAL ENCOUNTER|OBTURATOR SUBLUXATION OF UNSPECIFIED HIP, INITIAL ENCOUNTER
C2874008|T047|E09.638|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH OTHER ORAL COMPLICATIONS|DRUG/CHEM DIABETES MELLITUS W OTH ORAL COMPLICATIONS
C2833883|T037|S14.111D|ICD10CM|COMPLETE LESION AT C1 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION AT C1 LEVEL OF CERVICAL SPINAL CORD, SUBS
C2905674|T037|X72.XXXS|ICD10CM|INTENTIONAL SELF-HARM BY HANDGUN DISCHARGE, SEQUELA|INTENTIONAL SELF-HARM BY HANDGUN DISCHARGE, SEQUELA
C4269340|T037|S02.30XS|ICD10CM|FRACTURE OF ORBITAL FLOOR, UNSPECIFIED SIDE, SEQUELA|FRACTURE OF ORBITAL FLOOR, UNSPECIFIED SIDE, SEQUELA
C2901895|T047|M86.522|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, LEFT HUMERUS|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, LEFT HUMERUS
C2833882|T037|S14.111A|ICD10CM|COMPLETE LESION AT C1 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION AT C1 LEVEL OF CERVICAL SPINAL CORD, INIT
C4269468|T037|S02.621A|ICD10CM|FRACTURE OF SUBCONDYLAR PROCESS OF RIGHT MANDIBLE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF SUBCONDYLAR PROCESS OF RIGHT MANDIBLE, INIT
C2889577|T047|M08.419|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED SHOULDER|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED SHOULDER
C4269469|T037|S02.621B|ICD10CM|FRACTURE OF SUBCONDYLAR PROCESS OF RIGHT MANDIBLE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF SUBCONDYLAR PROCESS OF RIGHT MANDIBLE, 7THB
C2889576|T047|M08.412|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, LEFT SHOULDER|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, LEFT SHOULDER
C2889575|T047|M08.411|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, RIGHT SHOULDER|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, RIGHT SHOULDER
C2885205|T037|T61.92XA|ICD10CM|TOXIC EFFECT OF UNSPECIFIED SEAFOOD, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF UNSP SEAFOOD, INTENTIONAL SELF-HARM, INIT
C3264137|T033|Z89.512|ICD10CM|ACQUIRED ABSENCE OF LEFT LEG BELOW KNEE|ACQUIRED ABSENCE OF LEFT LEG BELOW KNEE
C2857993|T037|S72.345A|ICD10CM|NONDISPLACED SPIRAL FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED SPIRAL FRACTURE OF SHAFT OF LEFT FEMUR, INIT
C2857995|T037|S72.345C|ICD10CM|NONDISPLACED SPIRAL FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP SPIRAL FX SHAFT OF L FEMR, 7THC
C2857994|T037|S72.345B|ICD10CM|NONDISPLACED SPIRAL FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP SPIRAL FX SHAFT OF L FEMUR, INIT FOR OPN FX TYPE I/2
C2845984|T191|C7B.09|ICD10CM|SECONDARY CARCINOID TUMORS OF OTHER SITES|SECONDARY CARCINOID TUMORS OF OTHER SITES
C2845983|T191||ICD10CM|SECONDARY CARCINOID TUMORS OF PERITONEUM
C2845980|T191||ICD10CM|SECONDARY CARCINOID TUMORS OF DISTANT LYMPH NODES
C2845978|T191|C7B.00|ICD10CM|SECONDARY CARCINOID TUMORS, UNSPECIFIED SITE|SECONDARY CARCINOID TUMORS, UNSPECIFIED SITE
C2845982|T191||ICD10CM|SECONDARY CARCINOID TUMORS OF BONE
C2845981|T191||ICD10CM|SECONDARY CARCINOID TUMORS OF LIVER
C2901987|T046|M87.112|ICD10CM|OSTEONECROSIS DUE TO DRUGS, LEFT SHOULDER|OSTEONECROSIS DUE TO DRUGS, LEFT SHOULDER
C2911497|T033|Z94.84|ICD10CM|STEM CELLS TRANSPLANT STATUS|STEM CELLS TRANSPLANT STATUS
C2885339|T037|T63.022A|ICD10CM|TOXIC EFFECT OF CORAL SNAKE VENOM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CORAL SNAKE VENOM, SELF-HARM, INIT
C2911494|T033|Z94.81|ICD10CM|BONE MARROW TRANSPLANT STATUS|BONE MARROW TRANSPLANT STATUS
C2911495|T033|Z94.82|ICD10CM|INTESTINE TRANSPLANT STATUS|INTESTINE TRANSPLANT STATUS
C2911496|T033|Z94.83|ICD10CM|PANCREAS TRANSPLANT STATUS|PANCREAS TRANSPLANT STATUS
C2874793|T048|F19.121|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE ABUSE WITH INTOXICATION DELIRIUM|OTH PSYCHOACTIVE SUBSTANCE ABUSE WITH INTOXICATION DELIRIUM
C0839938|T047|M86.10|ICD10AM|OTHER ACUTE OSTEOMYELITIS, UNSPECIFIED SITE|OTHER ACUTE OSTEOMYELITIS, MULTIPLE SITES
C4268618|T047|K55.029|ICD10CM|ACUTE INFARCTION OF SMALL INTESTINE, EXTENT UNSPECIFIED|ACUTE INFARCTION OF SMALL INTESTINE, EXTENT UNSPECIFIED
C2832563|T037|S06.813S|ICD10CM|INJURY OF RIGHT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, SEQUELA|INJ R INT CAROTID, INTCR W LOC OF 1-5 HRS 59 MIN, SEQUELA
C2837840|T037|S32.313B|ICD10CM|DISPLACED AVULSION FRACTURE OF UNSPECIFIED ILIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISPLACED AVULSION FRACTURE OF UNSP ILIUM, INIT FOR OPN FX
C2889999|T037|T82.510A|ICD10CM|BREAKDOWN (MECHANICAL) OF SURGICALLY CREATED ARTERIOVENOUS FISTULA, INITIAL ENCOUNTER|BREAKDOWN OF SURGICALLY CREATED AV FISTULA, INIT
C2835378|T037|S22.061B|ICD10CM|STABLE BURST FRACTURE OF T7-T8 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|STABLE BURST FRACTURE OF T7-T8 VERTEBRA, INIT FOR OPN FX
C2890333|T037|T83.410A|ICD10CM|BREAKDOWN (MECHANICAL) OF IMPLANTED PENILE PROSTHESIS, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF IMPLANTED PENILE PROSTHESIS, INIT
C4268617|T047||ICD10CM|DIFFUSE ACUTE INFARCTION OF SMALL INTESTINE
C4268616|T047|K55.021|ICD10CM|FOCAL (SEGMENTAL) ACUTE INFARCTION OF SMALL INTESTINE|FOCAL (SEGMENTAL) ACUTE INFARCTION OF SMALL INTESTINE
C0392331|T048|F40.210|ICD10CM|ARACHNOPHOBIA|ARACHNOPHOBIA
C2874937|T048|F40.218|ICD10CM|OTHER ANIMAL TYPE PHOBIA|OTHER ANIMAL TYPE PHOBIA
C2835807|T037|S24.133S|ICD10CM|ANTERIOR CORD SYNDROME AT T7-T10 LEVEL OF THORACIC SPINAL CORD, SEQUELA|ANTERIOR CORD SYNDROME AT T7-T10, SEQUELA
C2858408|T037|S72.415C|ICD10CM|NONDISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP UNSP CONDYLE FX LOW END L FEMR, 7THC
C2901988|T046|M87.119|ICD10CM|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED SHOULDER|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED SHOULDER
C0085253|T047|M06.1|DMDICD10|ADULT-ONSET STILL'S DISEASE|ADULTE FORM DER STILL-KRANKHEIT
C2884184|T037|T52.92XA|ICD10CM|TOXIC EFFECT OF UNSPECIFIED ORGANIC SOLVENT, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF UNSP ORGANIC SOLVENT, SELF-HARM, INIT
C2890449|T037|T84.029A|ICD10CM|DISLOCATION OF UNSPECIFIED INTERNAL JOINT PROSTHESIS, INITIAL ENCOUNTER|DISLOCATION OF UNSP INTERNAL JOINT PROSTHESIS, INIT ENCNTR
C2834025|T037|S14.149A|ICD10CM|BROWN-SEQUARD SYNDROME AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|BROWN-SEQUARD SYND AT UNSP LEVEL OF CERV SPINAL CORD, INIT
C2884186|T037|T52.92XS|ICD10CM|TOXIC EFFECT OF UNSPECIFIED ORGANIC SOLVENT, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF UNSP ORGANIC SOLVENT, SELF-HARM, SEQUELA
C4268234|T048|F14.188|ICD10CM|COCAINE ABUSE WITH OTHER COCAINE-INDUCED DISORDER|COCAINE USE DISORDER, MILD, WITH COCAINE-INDUCED OBSESSIVE COMPULSIVE OR RELATED DISORDER
C4509284|T047|L97.205|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED CALF WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULCER OF UNSP CALF WITH MSL INVL W/O EVD OF NECR
C4509285|T047|L97.206|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED CALF WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OF UNSP CALF WITH BONE INVL W/O EVD OF NECR
C0348375|T191|C70|DMDICD10|MALIGNANT NEOPLASM OF MENINGES, UNSPECIFIED|BOESARTIGE NEUBILDUNG DER MENINGEN
C2832331|T037|S06.366S|ICD10CM|TRAUMATIC HEMORRHAGE OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|TRAUM HEMOR CEREB, W LOC >24 HR W/O RET CONSC W SURV, SQLA
C2888658|T047|L97.201|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED CALF LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHRONIC ULCER OF UNSP CALF LIMITED TO BRKDWN SKIN
C2888659|T047|L97.202|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED CALF WITH FAT LAYER EXPOSED|NON-PRESSURE CHRONIC ULCER OF UNSP CALF W FAT LAYER EXPOSED
C2888660|T047|L97.203|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED CALF WITH NECROSIS OF MUSCLE|NON-PRESSURE CHRONIC ULCER OF UNSP CALF W NECROSIS OF MUSCLE
C2874585|T048|F14.180|ICD10CM|COCAINE ABUSE WITH COCAINE-INDUCED ANXIETY DISORDER|COCAINE ABUSE WITH COCAINE-INDUCED ANXIETY DISORDER
C2874586|T048|F14.181|ICD10CM|COCAINE ABUSE WITH COCAINE-INDUCED SEXUAL DYSFUNCTION|COCAINE ABUSE WITH COCAINE-INDUCED SEXUAL DYSFUNCTION
C2874587|T048|F14.182|ICD10CM|COCAINE ABUSE WITH COCAINE-INDUCED SLEEP DISORDER|COCAINE ABUSE WITH COCAINE-INDUCED SLEEP DISORDER
C0153647|T191|C70.1|DMDICD10|MALIGNANT NEOPLASM OF SPINAL MENINGES|BOESARTIGE NEUBILDUNG: RUECKENMARKHAEUTE
C4509286|T047|L97.208|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED CALF WITH OTHER SPECIFIED SEVERITY|NON-PRS CHRONIC ULCER OF UNSPECIFIED CALF WITH OTH SEVERITY
C2888662|T047|L97.209|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED CALF WITH UNSPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF UNSP CALF WITH UNSP SEVERITY
C2877895|T037|T41.1X2S|ICD10CM|POISONING BY INTRAVENOUS ANESTHETICS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY INTRAVENOUS ANESTHETICS, SELF-HARM, SEQUELA
C2875080|T047|G40.019|ICD10CM|LOCALIZATION-RELATED (FOCAL) (PARTIAL) IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SEIZURES OF LOCALIZED ONSET, INTRACTABLE, WITHOUT STATUS EPILEPTICUS|LOCAL-REL IDIO EPI W SEIZ OF LOC ONSET, NTRCT, W/O STAT EPI
C2832105|T037|S06.312S|ICD10CM|CONTUSION AND LACERATION OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|CONTUS/LAC RIGHT CEREBRUM W LOC OF 31-59 MIN, SEQUELA
C2875079|T047|G40.011|ICD10CM|LOCALIZATION-RELATED (FOCAL) (PARTIAL) IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SEIZURES OF LOCALIZED ONSET, INTRACTABLE, WITH STATUS EPILEPTICUS|LOCAL-REL IDIO EPI W SEIZ OF LOC ONSET, NTRCT, W STAT EPI
C2890604|T037|T84.116A|ICD10CM|BREAKDOWN (MECHANICAL) OF INTERNAL FIXATION DEVICE OF BONE OF RIGHT LOWER LEG, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF INT FIX OF BONE OF R LOW LEG, INIT
C2889076|T047|M02.379|ICD10CM|REITER'S DISEASE, UNSPECIFIED ANKLE AND FOOT|REITER'S DISEASE, UNSPECIFIED ANKLE AND FOOT
C2835205|T037|S22.012B|ICD10CM|UNSTABLE BURST FRACTURE OF FIRST THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSTABLE BURST FX FIRST THOR VERTEBRA, INIT FOR OPN FX
C2835204|T037|S22.012A|ICD10CM|UNSTABLE BURST FRACTURE OF FIRST THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSTABLE BURST FRACTURE OF FIRST THORACIC VERTEBRA, INIT
C2874136|T047|E13.319|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH UNSPECIFIED DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA|OTH DIABETES W UNSP DIABETIC RETINOPATHY W/O MACULAR EDEMA
C0085222|T047|K68.12|ICD10CM|PSOAS MUSCLE ABSCESS|PSOAS MUSCLE ABSCESS
C2895206|T047|M35.9|ICD10CM|SYSTEMIC INVOLVEMENT OF CONNECTIVE TISSUE, UNSPECIFIED|AUTOIMMUNE DISEASE (SYSTEMIC) NOS
C0494951|T047|M35.8|DMDICD10|OTHER SPECIFIED SYSTEMIC INVOLVEMENT OF CONNECTIVE TISSUE|SONSTIGE NAEHER BEZEICHNETE KRANKHEITEN MIT SYSTEMBETEILIGUNG DES BINDEGEWEBES
C2889074|T047|M02.371|ICD10CM|REITER'S DISEASE, RIGHT ANKLE AND FOOT|REITER'S DISEASE, RIGHT ANKLE AND FOOT
C2883659|T037|T50.5X2A|ICD10CM|POISONING BY APPETITE DEPRESSANTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY APPETITE DEPRESSANTS, SELF-HARM, INIT
C0494949|T047|M35.5|DMDICD10|MULTIFOCAL FIBROSCLEROSIS|MULTIFOKALE FIBROSKLEROSE
C2889075|T047|M02.372|ICD10CM|REITER'S DISEASE, LEFT ANKLE AND FOOT|REITER'S DISEASE, LEFT ANKLE AND FOOT
C2874135|T047|E13.311|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH UNSPECIFIED DIABETIC RETINOPATHY WITH MACULAR EDEMA|OTH DIABETES W UNSP DIABETIC RETINOPATHY W MACULAR EDEMA
C0004943|T047|M35.2|DMDICD10|BEHCET'S DISEASE|BEHCET-KRANKHEIT
C1561633|T046|K68.19|ICD10CM|OTHER RETROPERITONEAL ABSCESS|OTHER RETROPERITONEAL ABSCESS
C2905662|T037|X71.8XXA|ICD10CM|OTHER INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION, INITIAL ENCOUNTER|OTH INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION, INIT
C2858165|T037|S72.363A|ICD10CM|DISPLACED SEGMENTAL FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED SEGMENTAL FRACTURE OF SHAFT OF UNSP FEMUR, INIT
C2858167|T037|S72.363C|ICD10CM|DISPLACED SEGMENTAL FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL SEG FX SHAFT OF UNSP FEMR, INIT FOR OPN FX TYPE 3A/B/C
C2858166|T037|S72.363B|ICD10CM|DISPLACED SEGMENTAL FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL SEG FX SHAFT OF UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2865530|T037|S88.021D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT KNEE LEVEL, RIGHT LOWER LEG, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION AT KNEE LEVEL, R LOW LEG, SUBS
C2832196|T037|S06.334S|ICD10CM|CONTUSION AND LACERATION OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|CONTUS/LAC CEREB, W LOC OF 6 HOURS TO 24 HOURS, SEQUELA
C2896552|T046|M80.041A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, RIGHT HAND, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, RIGHT HAND, INIT
C2845952|T191|C76.41|ICD10CM|MALIGNANT NEOPLASM OF RIGHT UPPER LIMB|MALIGNANT NEOPLASM OF RIGHT UPPER LIMB
C2845951|T191|C76.40|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED UPPER LIMB|MALIGNANT NEOPLASM OF UNSPECIFIED UPPER LIMB
C2845953|T191|C76.42|ICD10CM|MALIGNANT NEOPLASM OF LEFT UPPER LIMB|MALIGNANT NEOPLASM OF LEFT UPPER LIMB
C2902961|T047|N26.2|ICD10CM|PAGE KIDNEY|PAGE KIDNEY
C2838273|T037|S32.472B|ICD10CM|DISPLACED FRACTURE OF MEDIAL WALL OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISP FX OF MEDIAL WALL OF LEFT ACETABULUM, INIT FOR OPN FX
C2887185|T047|I83.015|ICD10CM|VARICOSE VEINS OF RIGHT LOWER EXTREMITY WITH ULCER OTHER PART OF FOOT|VARICOSE VEINS OF R LOW EXTREM W ULCER OTH PART OF FOOT
C2887183|T047|I83.014|ICD10CM|VARICOSE VEINS OF RIGHT LOWER EXTREMITY WITH ULCER OF HEEL AND MIDFOOT|VARICOSE VEINS OF R LOW EXTREM W ULCER OF HEEL AND MIDFOOT
C2887181|T047|I83.013|ICD10CM|VARICOSE VEINS OF RIGHT LOWER EXTREMITY WITH ULCER OF ANKLE|VARICOSE VEINS OF RIGHT LOWER EXTREMITY WITH ULCER OF ANKLE
C2887180|T047|I83.012|ICD10CM|VARICOSE VEINS OF RIGHT LOWER EXTREMITY WITH ULCER OF CALF|VARICOSE VEINS OF RIGHT LOWER EXTREMITY WITH ULCER OF CALF
C2887179|T047|I83.011|ICD10CM|VARICOSE VEINS OF RIGHT LOWER EXTREMITY WITH ULCER OF THIGH|VARICOSE VEINS OF RIGHT LOWER EXTREMITY WITH ULCER OF THIGH
C2860208|T037|S79.141A|ICD10CM|SALTER-HARRIS TYPE IV PHYSEAL FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SLTR-HARIS TYPE IV PHYSEAL FX LOWER END OF RIGHT FEMUR, INIT
C2887187|T047|I83.019|ICD10CM|VARICOSE VEINS OF RIGHT LOWER EXTREMITY WITH ULCER OF UNSPECIFIED SITE|VARICOSE VEINS OF RIGHT LOWER EXTREMITY W ULCER OF UNSP SITE
C2887186|T047|I83.018|ICD10CM|VARICOSE VEINS OF RIGHT LOWER EXTREMITY WITH ULCER OTHER PART OF LOWER LEG|VARICOSE VEINS OF R LOW EXTREM W ULCER OTH PART OF LOWER LEG
C2910356|T019|Q92.0|ICD10CM|WHOLE CHROMOSOME TRISOMY, NONMOSAICISM (MEIOTIC NONDISJUNCTION)|WHOLE CHROMOSOME TRISOMY, NONMOSAIC (MEIOTIC NONDISJUNCTION)
C2874121|T047||ICD10CM|TYPE 2 DIABETES MELLITUS WITH HYPOGLYCEMIA WITH COMA
C0348392|T191|C96.Z|ICD10CM|OTHER SPECIFIED MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE|OTH MALIG NEOPLM OF LYMPHOID, HEMATPOETC AND RELATED TISSUE
C2835760|T037|S24.102A|ICD10CM|UNSPECIFIED INJURY AT T2-T6 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY AT T2-T6 LEVEL OF THORACIC SPINAL CORD, INIT
C2832217|T037|S06.339S|ICD10CM|CONTUSION AND LACERATION OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|CONTUS/LAC CEREB, W LOC OF UNSP DURATION, SEQUELA
C4268276|T048|F18.17|ICD10CM|INHALANT ABUSE WITH INHALANT-INDUCED DEMENTIA|INHALANT USE DISORDER, MILD, WITH INHALANT INDUCED MAJOR NEUROCOGNITIVE DISORDER
C2905773|T037|X80.XXXA|ICD10CM|INTENTIONAL SELF-HARM BY JUMPING FROM A HIGH PLACE, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY JUMPING FROM A HIGH PLACE, INIT
C0334663|T191|C96.A|ICD10CM|HISTIOCYTIC SARCOMA|HISTIOCYTIC SARCOMA
C2874758|T048|F18.19|ICD10CM|INHALANT ABUSE WITH UNSPECIFIED INHALANT-INDUCED DISORDER|INHALANT ABUSE WITH UNSPECIFIED INHALANT-INDUCED DISORDER
C2896654|T046|M80.80XA|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, UNSPECIFIED SITE, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, UNSP SITE, INIT
C0027868|T047|G70.9|DMDICD10|MYONEURAL DISORDER, UNSPECIFIED|NEUROMUSKULAERE KRANKHEIT, NICHT NAEHER BEZEICHNET
C2861653|T191|C96.6|ICD10CM|UNIFOCAL LANGERHANS-CELL HISTIOCYTOSIS|HISTIOCYTOSIS X, UNIFOCAL
C2861650|T191|C96.4|ICD10CM|SARCOMA OF DENDRITIC CELLS (ACCESSORY CELLS)|SARCOMA OF DENDRITIC CELLS (ACCESSORY CELLS)
C2861652|T191|C96.5|ICD10CM|MULTIFOCAL AND UNISYSTEMIC LANGERHANS-CELL HISTIOCYTOSIS|MULTIFOCAL AND UNISYSTEMIC LANGERHANS-CELL HISTIOCYTOSIS
C0036221|T191|C96.2|DMDICD10|MALIGNANT MAST CELL TUMOR|BOESARTIGER MASTZELLTUMOR
C0268123|T047|E79.2|ICD10CM|MYOADENYLATE DEAMINASE DEFICIENCY|MYOADENYLATE DEAMINASE DEFICIENCY
C2861649|T191|C96.0|ICD10CM|MULTIFOCAL AND MULTISYSTEMIC (DISSEMINATED) LANGERHANS-CELL HISTIOCYTOSIS|MULTIFOCAL AND MULTISYSTEMIC LANGERHANS-CELL HISTIOCYTOSIS
C2893644|T047|M12.051|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], RIGHT HIP|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], RIGHT HIP
C2893645|T047|M12.052|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], LEFT HIP|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], LEFT HIP
C0034139|T047|E79|DMDICD10|DISORDER OF PURINE AND PYRIMIDINE METABOLISM, UNSPECIFIED|STOERUNGEN DES PURIN- UND PYRIMIDINSTOFFWECHSELS
C0348393|T191|C96.9|DMDICD10|MALIGNANT NEOPLASM OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE, UNSPECIFIED|BOESARTIGE NEUBILDUNG DES LYMPHATISCHEN, BLUTBILDENDEN UND VERWANDTEN GEWEBES, NICHT NAEHER BEZEICHNET
C2910366|T033|Q92.8|ICD10CM|OTHER SPECIFIED TRISOMIES AND PARTIAL TRISOMIES OF AUTOSOMES|DUPLICATIONS IDENTIFIED BY IN SITU HYBRIDIZATION (ISH)
C2838201|T037|S32.454B|ICD10CM|NONDISPLACED TRANSVERSE FRACTURE OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP TRANSVERSE FX RIGHT ACETABULUM, INIT FOR OPN FX
C2838200|T037|S32.454A|ICD10CM|NONDISPLACED TRANSVERSE FRACTURE OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED TRANSVERSE FRACTURE OF RIGHT ACETABULUM, INIT
C2837574|T037|S32.038A|ICD10CM|OTHER FRACTURE OF THIRD LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF THIRD LUMBAR VERTEBRA, INIT FOR CLOS FX
C2837575|T037|S32.038B|ICD10CM|OTHER FRACTURE OF THIRD LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF THIRD LUMBAR VERTEBRA, INIT FOR OPN FX
C0477675|T047|M83.5|DMDICD10|OTHER DRUG-INDUCED OSTEOMALACIA IN ADULTS|SONSTIGE ARZNEIMITTELINDUZIERTE OSTEOMALAZIE BEI ERWACHSENEN
C1442915|T047|K22.4|ICD10CM|DYSKINESIA OF ESOPHAGUS|CORKSCREW ESOPHAGUS
C2900587|T046|M83.2|ICD10CM|ADULT OSTEOMALACIA DUE TO MALABSORPTION|POSTSURGICAL MALABSORPTION OSTEOMALACIA IN ADULTS
C0451876|T047|M83.3|DMDICD10|ADULT OSTEOMALACIA DUE TO MALNUTRITION|OSTEOMALAZIE IM ERWACHSENENALTER DURCH FEHL- ODER MANGELERNAEHRUNG
C2900533|T046|M80.862A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, LEFT LOWER LEG, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, L LOW LEG, INIT
C2860156|T037|S79.119A|ICD10CM|SALTER-HARRIS TYPE I PHYSEAL FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SLTR-HARIS TYPE I PHYSEAL FX LOWER END OF UNSP FEMUR, INIT
C0686595|T191||ICD10AM|MONOCYTIC LEUKEMIA, UNSPECIFIED IN REMISSION
C2861625|T191|C93.90|ICD10CM|MONOCYTIC LEUKEMIA, UNSPECIFIED, NOT HAVING ACHIEVED REMISSION|MONOCYTIC LEUKEMIA, UNSP, NOT HAVING ACHIEVED REMISSION
C2349295|T191|C93.92|ICD10CM|MONOCYTIC LEUKEMIA, UNSPECIFIED IN RELAPSE|MONOCYTIC LEUKEMIA, UNSPECIFIED IN RELAPSE
C2882708|T047|I70.229|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES WITH REST PAIN, UNSPECIFIED EXTREMITY|ATHSCL NATIVE ARTERIES OF EXTRM W REST PAIN, UNSP EXTREMITY
C2879823|T037|T47.6X2S|ICD10CM|POISONING BY ANTIDIARRHEAL DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ANTIDIARRHEAL DRUGS, SELF-HARM, SEQUELA
C2874336|T048|F04|ICD10CM|AMNESTIC DISORDER DUE TO KNOWN PHYSIOLOGICAL CONDITION|AMNESTIC DISORDER DUE TO KNOWN PHYSIOLOGICAL CONDITION
C2888545|T047|L89.609|ICD10CM|PRESSURE ULCER OF UNSPECIFIED HEEL, UNSPECIFIED STAGE|PRESSURE ULCER OF UNSPECIFIED HEEL, UNSPECIFIED STAGE
C0153465|T191|C48.0|DMDICD10|MALIGNANT NEOPLASM OF RETROPERITONEUM|BOESARTIGE NEUBILDUNG: RETROPERITONEUM
C2888542|T047|L89.604|ICD10CM|PRESSURE ULCER OF UNSPECIFIED HEEL, STAGE 4|PRESSURE ULCER OF UNSPECIFIED HEEL, STAGE 4
C2349272|T191|C91.Z2|ICD10CM|OTHER LYMPHOID LEUKEMIA, IN RELAPSE|OTHER LYMPHOID LEUKEMIA, IN RELAPSE
C2888536|T047|L89.602|ICD10CM|PRESSURE ULCER OF UNSPECIFIED HEEL, STAGE 2|PRESSURE ULCER OF UNSPECIFIED HEEL, STAGE 2
C2854119|T191|C91.Z0|ICD10CM|OTHER LYMPHOID LEUKEMIA NOT HAVING ACHIEVED REMISSION|OTHER LYMPHOID LEUKEMIA NOT HAVING ACHIEVED REMISSION
C0153882|T191|C91.Z1|ICD10CM|OTHER LYMPHOID LEUKEMIA, IN REMISSION|OTHER LYMPHOID LEUKEMIA, IN REMISSION
C2945570|T033|Z99.2|DMDICD10|DEPENDENCE ON RENAL DIALYSIS|ABHAENGIGKEIT VON DIALYSE BEI NIERENINSUFFIZIENZ
C2882161|T047|I25.10|ICD10CM|ATHEROSCLEROTIC HEART DISEASE OF NATIVE CORONARY ARTERY WITHOUT ANGINA PECTORIS|ATHSCL HEART DISEASE OF NATIVE CORONARY ARTERY W/O ANG PCTRS
C2865550|T037|S88.119A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, UNSPECIFIED LOWER LEG, INITIAL ENCOUNTER|COMPLETE TRAUM AMP AT LEV BETW KN & ANKL, UNSP LOW LEG, INIT
C0006413|T191|C83.70|ICD10CM|BURKITT LYMPHOMA, UNSPECIFIED SITE|BURKITT LYMPHOMA, UNSPECIFIED SITE
C0153712|T191||ICD10CM|BURKITT LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK
C0153713|T191||ICD10CM|BURKITT LYMPHOMA, INTRATHORACIC LYMPH NODES
C0153714|T191||ICD10CM|BURKITT LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES
C0153715|T191||ICD10CM|BURKITT LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB
C0153716|T191|C83.75|ICD10CM|BURKITT LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|BURKITT LYMPHOMA, NODES OF INGUINAL REGION AND LOWER LIMB
C0153717|T191||ICD10CM|BURKITT LYMPHOMA, INTRAPELVIC LYMPH NODES
C0686546|T191||ICD10CM|BURKITT LYMPHOMA, SPLEEN
C0153719|T191||ICD10CM|BURKITT LYMPHOMA, LYMPH NODES OF MULTIPLE SITES
C2853932|T191||ICD10CM|BURKITT LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES
C2882704|T047|I70.221|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES WITH REST PAIN, RIGHT LEG|ATHSCL NATIVE ARTERIES OF EXTREMITIES W REST PAIN, RIGHT LEG
C2854080|T191||ICD10CM|EXTRAMEDULLARY PLASMACYTOMA IN RELAPSE
C0836956|T191||ICD10CM|EXTRAMEDULLARY PLASMACYTOMA IN REMISSION
C2854079|T191||ICD10CM|EXTRAMEDULLARY PLASMACYTOMA NOT HAVING ACHIEVED REMISSION
C2874133|T047|E13.29|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH OTHER DIABETIC KIDNEY COMPLICATION|OTH DIABETES MELLITUS WITH OTH DIABETIC KIDNEY COMPLICATION
C2865524|T037|S88.019A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT KNEE LEVEL, UNSPECIFIED LOWER LEG, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMP AT KNEE LEVEL, UNSP LOWER LEG, INIT
C2874131|T047|E13.22|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC CHRONIC KIDNEY DISEASE|OTH DIABETES MELLITUS WITH DIABETIC CHRONIC KIDNEY DISEASE
C2865525|T037|S88.019D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT KNEE LEVEL, UNSPECIFIED LOWER LEG, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMP AT KNEE LEVEL, UNSP LOWER LEG, SUBS
C2874130|T047|E13.21|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC NEPHROPATHY|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC NEPHROPATHY
C2865526|T037|S88.019S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT KNEE LEVEL, UNSPECIFIED LOWER LEG, SEQUELA|COMPLETE TRAUMATIC AMP AT KNEE LEVEL, UNSP LOW LEG, SEQUELA
C2858182|T037|S72.364A|ICD10CM|NONDISPLACED SEGMENTAL FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP SEGMENTAL FRACTURE OF SHAFT OF RIGHT FEMUR, INIT
C2910369|T049|Q93.7|ICD10CM|DELETIONS WITH OTHER COMPLEX REARRANGEMENTS|DELETIONS DUE TO UNBALANCED TRANSLOCATIONS, INVERSIONS AND INSERTIONS
C2875139|T047|G40.901|ICD10CM|EPILEPSY, UNSPECIFIED, NOT INTRACTABLE, WITH STATUS EPILEPTICUS|EPILEPSY, UNSP, NOT INTRACTABLE, WITH STATUS EPILEPTICUS
C2875140|T047|G40.909|ICD10CM|EPILEPSY, UNSPECIFIED, NOT INTRACTABLE, WITHOUT STATUS EPILEPTICUS|EPILEPSY, UNSP, NOT INTRACTABLE, WITHOUT STATUS EPILEPTICUS
C2879154|T037|T45.512S|ICD10CM|POISONING BY ANTICOAGULANTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ANTICOAGULANTS, INTENTIONAL SELF-HARM, SEQUELA
C0154408|T048||ICD10CM|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE, IN FULL REMISSION
C2874102|T047|E11.49|ICD10CM|TYPE 2 DIABETES MELLITUS WITH OTHER DIABETIC NEUROLOGICAL COMPLICATION|TYPE 2 DIABETES W OTH DIABETIC NEUROLOGICAL COMPLICATION
C2874916|T048||ICD10CM|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE, SEVERE WITH PSYCHOTIC FEATURES
C0494399|T048|F32.2|DMDICD10|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE, SEVERE WITHOUT PSYCHOTIC FEATURES|SCHWERE DEPRESSIVE EPISODE OHNE PSYCHOTISCHE SYMPTOME
C0494398|T048|F32.1|DMDICD10|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE, MODERATE|MITTELGRADIGE DEPRESSIVE EPISODE
C2888319|T047|L89.134|ICD10CM|PRESSURE ULCER OF RIGHT LOWER BACK, STAGE 4|PRESSURE ULCER OF RIGHT LOWER BACK, STAGE 4
C2874098|T047|E11.42|ICD10CM|TYPE 2 DIABETES MELLITUS WITH DIABETIC POLYNEUROPATHY|TYPE 2 DIABETES MELLITUS WITH DIABETIC NEURALGIA
C2874100|T047|E11.43|ICD10CM|TYPE 2 DIABETES MELLITUS WITH DIABETIC AUTONOMIC (POLY)NEUROPATHY|TYPE 2 DIABETES W DIABETIC AUTONOMIC (POLY)NEUROPATHY
C2874097|T047|E11.40|ICD10CM|TYPE 2 DIABETES MELLITUS WITH DIABETIC NEUROPATHY, UNSPECIFIED|TYPE 2 DIABETES MELLITUS WITH DIABETIC NEUROPATHY, UNSP
C0837043|T047|E11.41|ICD10AM|TYPE 2 DIABETES MELLITUS WITH DIABETIC MONONEUROPATHY|TYPE 2 DIABETES MELLITUS WITH DIABETIC MONONEUROPATHY
C2883861|T037|T50.A92A|ICD10CM|POISONING BY OTHER BACTERIAL VACCINES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH BACTERIAL VACCINES, SELF-HARM, INIT
C1269683|T048||ICD10CM|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE, UNSPECIFIED
C2832586|T037|S06.819A|ICD10CM|INJURY OF RIGHT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|INJURY OF R INT CAROTID, INTCR W LOC OF UNSP DURATION, INIT
C2879152|T037|T45.512A|ICD10CM|POISONING BY ANTICOAGULANTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ANTICOAGULANTS, INTENTIONAL SELF-HARM, INIT
C2887903|T047|K63.1|ICD10CM|PERFORATION OF INTESTINE (NONTRAUMATIC)|PERFORATION (NONTRAUMATIC) OF RECTUM
C2884593|T037|T56.812A|ICD10CM|TOXIC EFFECT OF THALLIUM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF THALLIUM, INTENTIONAL SELF-HARM, INIT ENCNTR
C2883863|T037|T50.A92S|ICD10CM|POISONING BY OTHER BACTERIAL VACCINES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH BACTERIAL VACCINES, SELF-HARM, SEQUELA
C2882349|T047|I63.139|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF UNSPECIFIED CAROTID ARTERY|CEREBRAL INFARCTION DUE TO EMBOLISM OF UNSP CAROTID ARTERY
C2891319|T037|T87.0X2|ICD10CM|COMPLICATIONS OF REATTACHED (PART OF) LEFT UPPER EXTREMITY|COMPLICATIONS OF REATTACHED (PART OF) LEFT UPPER EXTREMITY
C2891318|T037|T87.0X1|ICD10CM|COMPLICATIONS OF REATTACHED (PART OF) RIGHT UPPER EXTREMITY|COMPLICATIONS OF REATTACHED (PART OF) RIGHT UPPER EXTREMITY
C3463824|T191|D46.9|DMDICD10|MYELODYSPLASTIC SYNDROME, UNSPECIFIED|MYELODYSPLASTISCHES SYNDROM, NICHT NAEHER BEZEICHNET
C2882348|T047|I63.132|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF LEFT CAROTID ARTERY|CEREBRAL INFARCTION DUE TO EMBOLISM OF LEFT CAROTID ARTERY
C4268478|T047|I63.133|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF BILATERAL CAROTID ARTERIES|CEREBRAL INFRC DUE TO EMBOLISM OF BILATERAL CAROTID ARTERIES
C0348439|T191|D46.4|DMDICD10|REFRACTORY ANEMIA, UNSPECIFIED|REFRAKTAERE ANAEMIE, NICHT NAEHER BEZEICHNET
C2882347|T047|I63.131|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF RIGHT CAROTID ARTERY|CEREBRAL INFARCTION DUE TO EMBOLISM OF RIGHT CAROTID ARTERY
C2873713|T191|D46.0|ICD10CM|REFRACTORY ANEMIA WITHOUT RING SIDEROBLASTS, SO STATED|REFRACTORY ANEMIA WITHOUT RING SIDEROBLASTS, SO STATED
C1264195|T191|D46.1|ICD10CM|REFRACTORY ANEMIA WITH RING SIDEROBLASTS|REFRACTORY ANEMIA WITH RING SIDEROBLASTS
C2842090|T191|C50.129|ICD10CM|MALIGNANT NEOPLASM OF CENTRAL PORTION OF UNSPECIFIED MALE BREAST|MALIGNANT NEOPLASM OF CENTRAL PORTION OF UNSP MALE BREAST
C3264197|T047|H40.1221|ICD10CM|LOW-TENSION GLAUCOMA, LEFT EYE, MILD STAGE|LOW-TENSION GLAUCOMA, LEFT EYE, MILD STAGE
C3264198|T047|H40.1222|ICD10CM|LOW-TENSION GLAUCOMA, LEFT EYE, MODERATE STAGE|LOW-TENSION GLAUCOMA, LEFT EYE, MODERATE STAGE
C3264199|T047|H40.1223|ICD10CM|LOW-TENSION GLAUCOMA, LEFT EYE, SEVERE STAGE|LOW-TENSION GLAUCOMA, LEFT EYE, SEVERE STAGE
C3264200|T047|H40.1224|ICD10CM|LOW-TENSION GLAUCOMA, LEFT EYE, INDETERMINATE STAGE|LOW-TENSION GLAUCOMA, LEFT EYE, INDETERMINATE STAGE
C2842088|T191|C50.121|ICD10CM|MALIGNANT NEOPLASM OF CENTRAL PORTION OF RIGHT MALE BREAST|MALIGNANT NEOPLASM OF CENTRAL PORTION OF RIGHT MALE BREAST
C2842089|T191|C50.122|ICD10CM|MALIGNANT NEOPLASM OF CENTRAL PORTION OF LEFT MALE BREAST|MALIGNANT NEOPLASM OF CENTRAL PORTION OF LEFT MALE BREAST
C2855907|T037|S68.120S|ICD10CM|PARTIAL TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF RIGHT INDEX FINGER, SEQUELA|PARTIAL TRAUMATIC MCP AMPUTATION OF R IDX FNGR, SEQUELA
C0010314|T047|Q93.4|DMDICD10|DELETION OF SHORT ARM OF CHROMOSOME 5|DELETION DES KURZEN ARMES DES CHROMOSOMS 5
C0494210|T191|D46.Z|ICD10CM|OTHER MYELODYSPLASTIC SYNDROMES|OTHER MYELODYSPLASTIC SYNDROMES
C2832616|T037|S06.826S|ICD10CM|INJURY OF LEFT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|INJ L INT CRTD,INTCR W LOC >24 HR W/O RET CONSC W SURV, SQLA
C2860244|T037|S79.199A|ICD10CM|OTHER PHYSEAL FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH PHYSEAL FRACTURE OF LOWER END OF UNSP FEMUR, INIT
C2882432|T047|I66.13|ICD10CM|OCCLUSION AND STENOSIS OF BILATERAL ANTERIOR CEREBRAL ARTERIES|OCCLUSION AND STENOSIS OF BI ANTERIOR CEREBRAL ARTERIES
C2882431|T047|I66.12|ICD10CM|OCCLUSION AND STENOSIS OF LEFT ANTERIOR CEREBRAL ARTERY|OCCLUSION AND STENOSIS OF LEFT ANTERIOR CEREBRAL ARTERY
C2882430|T047|I66.11|ICD10CM|OCCLUSION AND STENOSIS OF RIGHT ANTERIOR CEREBRAL ARTERY|OCCLUSION AND STENOSIS OF RIGHT ANTERIOR CEREBRAL ARTERY
C2853814|T191|C82.28|ICD10CM|FOLLICULAR LYMPHOMA GRADE III, UNSPECIFIED, LYMPH NODES OF MULTIPLE SITES|FOLLICULAR LYMPHOMA GRADE III, UNSP, LYMPH NODES MULT SITE
C2832614|T037|S06.826A|ICD10CM|INJURY OF LEFT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|INJ L INT CRTD,INTCR W LOC >24 HR W/O RET CONSC W SURV, INIT
C2874280|T047|E76.21|ICD10CM|MORQUIO MUCOPOLYSACCHARIDOSES, UNSPECIFIED|MORQUIO MUCOPOLYSACCHARIDOSES
C2882433|T047|I66.19|ICD10CM|OCCLUSION AND STENOSIS OF UNSPECIFIED ANTERIOR CEREBRAL ARTERY|OCCLUSION AND STENOSIS OF UNSP ANTERIOR CEREBRAL ARTERY
C2853815|T191|C82.29|ICD10CM|FOLLICULAR LYMPHOMA GRADE III, UNSPECIFIED, EXTRANODAL AND SOLID ORGAN SITES|FOLICLAR LYMPH GRADE III, UNSP, EXTRNOD AND SOLID ORG SITES
C1301356|T191|D46.B|ICD10CM|REFRACTORY CYTOPENIA WITH MULTILINEAGE DYSPLASIA AND RING SIDEROBLASTS|REFRACT CYTOPENIA W MULTILIN DYSPLASIA AND RING SIDEROBLASTS
C1292779|T191|D46.C|ICD10CM|MYELODYSPLASTIC SYNDROME WITH ISOLATED DEL(5Q) CHROMOSOMAL ABNORMALITY|MYELODYSPLASTIC SYNDROME W ISOLATED DEL(5Q) CHROMSOML ABNLT
C0796466|T191|D46.A|ICD10CM|REFRACTORY CYTOPENIA WITH MULTILINEAGE DYSPLASIA|REFRACTORY CYTOPENIA WITH MULTILINEAGE DYSPLASIA
C2889219|T047|M05.352|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT HIP|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF LEFT HIP
C2883133|T047|I82.539|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED POPLITEAL VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF UNSP POPLITEAL VEIN
C2889218|T047|M05.351|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT HIP|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF RIGHT HIP
C2883132|T047|I82.533|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF POPLITEAL VEIN, BILATERAL|CHRONIC EMBOLISM AND THROMBOSIS OF POPLITEAL VEIN, BILATERAL
C2883131|T047|I82.532|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF LEFT POPLITEAL VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF LEFT POPLITEAL VEIN
C2883130|T047|I82.531|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF RIGHT POPLITEAL VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF RIGHT POPLITEAL VEIN
C2889217|T047|M05.359|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP
C2856109|T037|S68.729S|ICD10CM|PARTIAL TRAUMATIC TRANSMETACARPAL AMPUTATION OF UNSPECIFIED HAND, SEQUELA|PARTIAL TRAUMATIC TRANSMETCRPL AMP OF UNSP HAND, SEQUELA
C2878330|T037|T43.1X2S|ICD10CM|POISONING BY MONOAMINE-OXIDASE-INHIBITOR ANTIDEPRESSANTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY MAO INHIB ANTIDEPRESSANTS, SELF-HARM, SEQUELA
C2876820|T037|T37.1X2S|ICD10CM|POISONING BY ANTIMYCOBACTERIAL DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ANTIMYCOBACTERIAL DRUGS, SELF-HARM, SEQUELA
C0016952|T047||ICD10CM|GALACTOSEMIA
C0342745|T047|E74.20|ICD10CM|DISORDERS OF GALACTOSE METABOLISM, UNSPECIFIED|DISORDERS OF GALACTOSE METABOLISM, UNSPECIFIED
C2874279|T047|E76.211|ICD10CM|MORQUIO B MUCOPOLYSACCHARIDOSES|MORQUIO B MUCOPOLYSACCHARIDOSES
C2874269|T047|E74.29|ICD10CM|OTHER DISORDERS OF GALACTOSE METABOLISM|OTHER DISORDERS OF GALACTOSE METABOLISM
C3263946|T047|D68.318|ICD10CM|OTHER HEMORRHAGIC DISORDER DUE TO INTRINSIC CIRCULATING ANTICOAGULANTS, ANTIBODIES, OR INHIBITORS|HEMORRHAGIC DISORDER DUE TO INTRINSIC INCREASE IN ANTITHROMBIN
C2882414|T047|I63.549|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF UNSPECIFIED CEREBELLAR ARTERY|CEREB INFRC DUE TO UNSP OCCLS OR STENOS OF UNSP CEREBLR ART
C4268492|T047|I63.543|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF BILATERAL CEREBELLAR ARTERIES|CEREB INFRC DUE TO UNSP OCCLS OR STENOSIS OF BI CEREBLR ART
C2882413|T047|I63.542|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF LEFT CEREBELLAR ARTERY|CEREB INFRC DUE TO UNSP OCCLS OR STENOS OF LEFT CEREBLR ART
C2882412|T047|I63.541|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF RIGHT CEREBELLAR ARTERY|CEREB INFRC DUE TO UNSP OCCLS OR STENOS OF RIGHT CEREBLR ART
C4269392|T037|S02.40CB|ICD10CM|MAXILLARY FRACTURE, RIGHT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|MAXILLARY FRACTURE, RIGHT SIDE, 7THB
C2873805|T047|D69.1|ICD10CM|QUALITATIVE PLATELET DEFECTS|THROMBOASTHENIA (HEMORRHAGIC) (HEREDITARY)
C2833339|T037|S12.231B|ICD10CM|UNSPECIFIED TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP TRAUM NONDISP SPONDYLOLYSIS OF 3RD CERVCAL VERT, 7THB
C0348836|T047|I66.3|DMDICD10|OCCLUSION AND STENOSIS OF CEREBELLAR ARTERIES|VERSCHLUSS UND STENOSE DER AA. CEREBELLI
C2875151|T047|G43.109|ICD10CM|MIGRAINE WITH AURA, NOT INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|MIGRAINE WITH AURA, NOT INTRACTABLE, W/O STATUS MIGRAINOSUS
C1368065|T046|D69.0|ICD10CM|ALLERGIC PURPURA|VASCULAR PURPURA
C2901103|T046|M84.477A|ICD10CM|PATHOLOGICAL FRACTURE, RIGHT TOE(S), INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, RIGHT TOE(S), INIT FOR FX
C2875150|T047|G43.101|ICD10CM|MIGRAINE WITH AURA, NOT INTRACTABLE, WITH STATUS MIGRAINOSUS|MIGRAINE WITH AURA, NOT INTRACTABLE, WITH STATUS MIGRAINOSUS
C2882438|T047|I66.8|ICD10CM|OCCLUSION AND STENOSIS OF OTHER CEREBRAL ARTERIES|OCCLUSION AND STENOSIS OF PERFORATING ARTERIES
C0272309|T047|D69.2|ICD10CM|OTHER NONTHROMBOCYTOPENIC PURPURA|PURPURA SIMPLEX
C0694509|T047|K87|DMDICD10|DISORDERS OF GALLBLADDER, BILIARY TRACT AND PANCREAS IN DISEASES CLASSIFIED ELSEWHERE|KRANKHEITEN DER GALLENBLASE, DER GALLENWEGE UND DES PANKREAS BEI ANDERENORTS KLASSIFIZIERTEN KRANKHEITEN
C2832669|T037|S06.899S|ICD10CM|OTHER SPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|INTCRAN INJ W LOC OF UNSP DURATION, SEQUELA
C2911501|T033|Z95.811|ICD10CM|PRESENCE OF HEART ASSIST DEVICE|PRESENCE OF HEART ASSIST DEVICE
C2885543|T037|T63.312S|ICD10CM|TOXIC EFFECT OF VENOM OF BLACK WIDOW SPIDER, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF BLACK WIDOW SPIDER, SLF-HRM, SQLA
C2911502|T033|Z95.812|ICD10CM|PRESENCE OF FULLY IMPLANTABLE ARTIFICIAL HEART|PRESENCE OF FULLY IMPLANTABLE ARTIFICIAL HEART
C0600433|T047||ICD10CM|ACTIVATED PROTEIN C RESISTANCE
C1260403|T047||ICD10CM|PROTHROMBIN GENE MUTATION
C2837817|T037|S32.309A|ICD10CM|UNSPECIFIED FRACTURE OF UNSPECIFIED ILIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF UNSP ILIUM, INIT ENCNTR FOR CLOSED FRACTURE
C2837818|T037|S32.309B|ICD10CM|UNSPECIFIED FRACTURE OF UNSPECIFIED ILIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF UNSP ILIUM, INIT ENCNTR FOR OPEN FRACTURE
C2873799|T046|D68.59|ICD10CM|OTHER PRIMARY THROMBOPHILIA|OTHER PRIMARY THROMBOPHILIA
C0494456|T047|G13.8|DMDICD10|SYSTEMIC ATROPHY PRIMARILY AFFECTING CENTRAL NERVOUS SYSTEM IN OTHER DISEASES CLASSIFIED ELSEWHERE|SYSTEMATROPHIEN, VORWIEGEND DAS ZENTRALNERVENSYSTEM BETREFFEND, BEI SONSTIGEN ANDERENORTS KLASSIFIZIERTEN KRANKHEITEN
C2882799|T047|I70.398|ICD10CM|OTHER ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, OTHER EXTREMITY|OTH ATHSCL UNSP TYPE BYPASS OF THE EXTRM, OTH EXTREMITY
C2882800|T047|I70.399|ICD10CM|OTHER ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, UNSPECIFIED EXTREMITY|OTH ATHSCL UNSP TYPE BYPASS OF THE EXTRM, UNSP EXTREMITY
C2875377|T047|G90.529|ICD10CM|COMPLEX REGIONAL PAIN SYNDROME I OF UNSPECIFIED LOWER LIMB|COMPLEX REGIONAL PAIN SYNDROME I OF UNSPECIFIED LOWER LIMB
C2911408|T033|Z89.419|ICD10CM|ACQUIRED ABSENCE OF UNSPECIFIED GREAT TOE|ACQUIRED ABSENCE OF UNSPECIFIED GREAT TOE
C2878305|T037|T43.022S|ICD10CM|POISONING BY TETRACYCLIC ANTIDEPRESSANTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY TETRACYCLIC ANTIDEPRESSANTS, SELF-HARM, SEQUELA
C0494454|T047|G13.1|DMDICD10|OTHER SYSTEMIC ATROPHY PRIMARILY AFFECTING CENTRAL NERVOUS SYSTEM IN NEOPLASTIC DISEASE|SONSTIGE SYSTEMATROPHIEN, VORWIEGEND DAS ZENTRALNERVENSYSTEM BETREFFEND, BEI NEUBILDUNGEN
C2875053|T047|G13.0|ICD10CM|PARANEOPLASTIC NEUROMYOPATHY AND NEUROPATHY|SENSORIAL PARANEOPLASTIC NEUROPATHY [DENNY BROWN]
C0494455|T047|G13.2|DMDICD10|SYSTEMIC ATROPHY PRIMARILY AFFECTING THE CENTRAL NERVOUS SYSTEM IN MYXEDEMA|SYSTEMATROPHIE, VORWIEGEND DAS ZENTRALNERVENSYSTEM BETREFFEND, BEI MYXOEDEM
C2875374|T047|G90.521|ICD10CM|COMPLEX REGIONAL PAIN SYNDROME I OF RIGHT LOWER LIMB|COMPLEX REGIONAL PAIN SYNDROME I OF RIGHT LOWER LIMB
C2911406|T033|Z89.411|ICD10CM|ACQUIRED ABSENCE OF RIGHT GREAT TOE|ACQUIRED ABSENCE OF RIGHT GREAT TOE
C2875376|T047|G90.523|ICD10CM|COMPLEX REGIONAL PAIN SYNDROME I OF LOWER LIMB, BILATERAL|COMPLEX REGIONAL PAIN SYNDROME I OF LOWER LIMB, BILATERAL
C2875375|T047|G90.522|ICD10CM|COMPLEX REGIONAL PAIN SYNDROME I OF LEFT LOWER LIMB|COMPLEX REGIONAL PAIN SYNDROME I OF LEFT LOWER LIMB
C2887788|T047|K51.00|ICD10CM|ULCERATIVE (CHRONIC) PANCOLITIS WITHOUT COMPLICATIONS|ULCERATIVE (CHRONIC) PANCOLITIS WITHOUT COMPLICATIONS
C2878303|T037|T43.022A|ICD10CM|POISONING BY TETRACYCLIC ANTIDEPRESSANTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY TETRACYCLIC ANTIDEPRESSANTS, SELF-HARM, INIT
C4269445|T037|S02.610S|ICD10CM|FRACTURE OF CONDYLAR PROCESS OF MANDIBLE, UNSPECIFIED SIDE, SEQUELA|FX CONDYLAR PROCESS OF MANDIBLE, UNSPECIFIED SIDE, SEQUELA
C4509207|T047|I27.0|ICD10CM|PRIMARY PULMONARY HYPERTENSION|PRIMARY PULMONARY ARTERIAL HYPERTENSION
C0152102|T047|I27.1|DMDICD10|KYPHOSCOLIOTIC HEART DISEASE|KYPHOSKOLIOTISCHE HERZKRANKHEIT
C2882223|T047|I27.29|ICD10CM|OTHER SECONDARY PULMONARY HYPERTENSION|OTHER SECONDARY PULMONARY HYPERTENSION
C4269441|T037|S02.610B|ICD10CM|FRACTURE OF CONDYLAR PROCESS OF MANDIBLE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FX CONDYLAR PROCESS OF MANDIBLE, UNSPECIFIED SIDE, 7THB
C2835457|T037|S22.082B|ICD10CM|UNSTABLE BURST FRACTURE OF T11-T12 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSTABLE BURST FRACTURE OF T11-T12 VERTEBRA, INIT FOR OPN FX
C2835456|T037|S22.082A|ICD10CM|UNSTABLE BURST FRACTURE OF T11-T12 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSTABLE BURST FRACTURE OF T11-T12 VERTEBRA, INIT
C0238074|T047|I27.9|ICD10CM|PULMONARY HEART DISEASE, UNSPECIFIED|CHRONIC CARDIOPULMONARY DISEASE
C2853890|T191|C83.06|ICD10CM|SMALL CELL B-CELL LYMPHOMA, INTRAPELVIC LYMPH NODES|SMALL CELL B-CELL LYMPHOMA, INTRAPELVIC LYMPH NODES
C0153506|T191|C39.0|DMDICD10|MALIGNANT NEOPLASM OF UPPER RESPIRATORY TRACT, PART UNSPECIFIED|BOESARTIGE NEUBILDUNG: OBERE ATEMWEGE, TEIL NICHT NAEHER BEZEICHNET
C0275583|T047|A43.0|DMDICD10|PULMONARY NOCARDIOSIS|PULMONALE NOKARDIOSE
C2886159|T037|T65.822A|ICD10CM|TOXIC EFFECT OF HARMFUL ALGAE AND ALGAE TOXINS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFF OF HARMFUL ALGAE AND ALGAE TOXINS, SLF-HRM, INIT
C2837964|T191|C39.9|ICD10CM|MALIGNANT NEOPLASM OF LOWER RESPIRATORY TRACT, PART UNSPECIFIED|MALIGNANT NEOPLASM OF LOWER RESPIRATORY TRACT, PART UNSP
C2875328|T184||ICD10CM|FLACCID HEMIPLEGIA AFFECTING RIGHT NONDOMINANT SIDE
C2875327|T184||ICD10CM|FLACCID HEMIPLEGIA AFFECTING LEFT DOMINANT SIDE
C2875326|T184||ICD10CM|FLACCID HEMIPLEGIA AFFECTING RIGHT DOMINANT SIDE
C0154693|T184|G81.00|ICD10CM|FLACCID HEMIPLEGIA AFFECTING UNSPECIFIED SIDE|FLACCID HEMIPLEGIA AFFECTING UNSPECIFIED SIDE
C2875329|T184||ICD10CM|FLACCID HEMIPLEGIA AFFECTING LEFT NONDOMINANT SIDE
C2905819|T037|X83.8XXS|ICD10CM|INTENTIONAL SELF-HARM BY OTHER SPECIFIED MEANS, SEQUELA|INTENTIONAL SELF-HARM BY OTHER SPECIFIED MEANS, SEQUELA
C2878482|T037|T43.4X2A|ICD10CM|POISONING BY BUTYROPHENONE AND THIOTHIXENE NEUROLEPTICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY BUTYROPHEN/THIOTHIXEN NEUROLEPTC, SELF-HARM, INIT
C2889410|T047|M06.072|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, LEFT ANKLE AND FOOT|RHEUMATOID ARTHRITIS W/O RHEUMATOID FACTOR, LEFT ANK/FT
C2887276|T047|I87.019|ICD10CM|POSTTHROMBOTIC SYNDROME WITH ULCER OF UNSPECIFIED LOWER EXTREMITY|POSTTHROMBOTIC SYNDROME WITH ULCER OF UNSP LOWER EXTREMITY
C2889409|T047|M06.071|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, RIGHT ANKLE AND FOOT|RHEUMATOID ARTHRITIS W/O RHEUMATOID FACTOR, RIGHT ANK/FT
C2887275|T047|I87.013|ICD10CM|POSTTHROMBOTIC SYNDROME WITH ULCER OF BILATERAL LOWER EXTREMITY|POSTTHROMBOTIC SYNDROME W ULCER OF BILATERAL LOWER EXTREMITY
C2887274|T047|I87.012|ICD10CM|POSTTHROMBOTIC SYNDROME WITH ULCER OF LEFT LOWER EXTREMITY|POSTTHROMBOTIC SYNDROME WITH ULCER OF LEFT LOWER EXTREMITY
C2887273|T047|I87.011|ICD10CM|POSTTHROMBOTIC SYNDROME WITH ULCER OF RIGHT LOWER EXTREMITY|POSTTHROMBOTIC SYNDROME WITH ULCER OF RIGHT LOWER EXTREMITY
C2889411|T047|M06.079|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, UNSPECIFIED ANKLE AND FOOT|RHEUMATOID ARTHRITIS W/O RHEUMATOID FACTOR, UNSP ANK/FT
C2890538|T037|T84.062A|ICD10CM|WEAR OF ARTICULAR BEARING SURFACE OF INTERNAL PROSTHETIC RIGHT KNEE JOINT, INITIAL ENCOUNTER|WEAR OF ARTIC BEARING SURFACE OF INT PROSTH R KNEE JT, INIT
C2890099|T037|T82.590A|ICD10CM|OTHER MECHANICAL COMPLICATION OF SURGICALLY CREATED ARTERIOVENOUS FISTULA, INITIAL ENCOUNTER|MECH COMPL OF SURGICALLY CREATED ARTERIOVENOUS FISTULA, INIT
C2896604|T046|M80.062A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, LEFT LOWER LEG, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, L LOW LEG, INIT
C2900867|T046|M84.411A|ICD10CM|PATHOLOGICAL FRACTURE, RIGHT SHOULDER, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, RIGHT SHOULDER, INIT FOR FX
C2874014|T047|E09.8|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH UNSPECIFIED COMPLICATIONS|DRUG/CHEM DIABETES MELLITUS W UNSP COMPLICATIONS
C2874015|T047|E09.9|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITHOUT COMPLICATIONS|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS W/O COMPLICATIONS
C0864959|T191|C57.9|ICD10CM|MALIGNANT NEOPLASM OF FEMALE GENITAL ORGAN, UNSPECIFIED|MALIGNANT NEOPLASM OF FEMALE GENITOURINARY TRACT NOS
C2842160|T191|C57.8|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF FEMALE GENITAL ORGANS|PRIMARY UTERO-OVARIAN MALIGNANT NEOPLASM WHOSE POINT OF ORIGIN CANNOT BE DETERMINED
C0153584|T191|C57.4|DMDICD10|MALIGNANT NEOPLASM OF UTERINE ADNEXA, UNSPECIFIED|BOESARTIGE NEUBILDUNG: UTERINE ADNEXE, NICHT NAEHER BEZEICHNET
C2842157|T191|C57.7|ICD10CM|MALIGNANT NEOPLASM OF OTHER SPECIFIED FEMALE GENITAL ORGANS|MALIGNANT NEOPLASM OF WOLFFIAN BODY OR DUCT
C0864950|T191||ICD10CM|MALIGNANT NEOPLASM OF PARAMETRIUM
C2830236|T047|B42.82|ICD10CM|SPOROTRICHOSIS ARTHRITIS|SPOROTRICHOSIS ARTHRITIS
C0600452|T047||ICD10CM|HEPATOPULMONARY SYNDROME
C2889973|T037|T82.399A|ICD10CM|OTHER MECHANICAL COMPLICATION OF UNSPECIFIED VASCULAR GRAFTS, INITIAL ENCOUNTER|MECH COMPL OF UNSPECIFIED VASCULAR GRAFTS, INITIAL ENCOUNTER
C2891324|T037|T87.30|ICD10CM|NEUROMA OF AMPUTATION STUMP, UNSPECIFIED EXTREMITY|NEUROMA OF AMPUTATION STUMP, UNSPECIFIED EXTREMITY
C2874315|T046|E89.0|ICD10CM|POSTPROCEDURAL HYPOTHYROIDISM|POSTIRRADIATION HYPOTHYROIDISM
C2832286|T037|S06.356A|ICD10CM|TRAUMATIC HEMORRHAGE OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|TRAUM HEMOR L CEREB W LOC >24 HR W/O RET CONSC W SURV, INIT
C2058370|T037||MTHICD9|POSTPROCEDURAL HYPOPARATHYROIDISM
C2874316|T046|E89.3|ICD10CM|POSTPROCEDURAL HYPOPITUITARISM|POSTIRRADIATION HYPOPITUITARISM
C3887666|T047|E32.0|DMDICD10|PERSISTENT HYPERPLASIA OF THYMUS|PERSISTIERENDE THYMUSHYPERPLASIE
C0154200|T047|E32.1|DMDICD10|ABSCESS OF THYMUS|ABSZESS DES THYMUS
C0348465|T047|E32.8|DMDICD10|OTHER DISEASES OF THYMUS|SONSTIGE KRANKHEITEN DES THYMUS
C0154199|T047|E32|DMDICD10|DISEASE OF THYMUS, UNSPECIFIED|KRANKHEITEN DES THYMUS
C2859988|T037|S78.022A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEFT HIP JOINT, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION AT LEFT HIP JOINT, INIT ENCNTR
C2876212|T037|T32.73|ICD10CM|CORROSIONS INVOLVING 70-79% OF BODY SURFACE WITH 30-39% THIRD DEGREE CORROSION|CORROS 70-79% OF BODY SURFACE W 30-39% THIRD DEGREE CORROS
C2832288|T037|S06.356S|ICD10CM|TRAUMATIC HEMORRHAGE OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|TRAUM HEMOR L CEREB W LOC >24 HR W/O RET CONSC W SURV, SQLA
C2859989|T037|S78.022D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEFT HIP JOINT, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION AT LEFT HIP JOINT, SUBS ENCNTR
C2876211|T037|T32.72|ICD10CM|CORROSIONS INVOLVING 70-79% OF BODY SURFACE WITH 20-29% THIRD DEGREE CORROSION|CORROS 70-79% OF BODY SURFACE W 20-29% THIRD DEGREE CORROS
C2876210|T037|T32.71|ICD10CM|CORROSIONS INVOLVING 70-79% OF BODY SURFACE WITH 10-19% THIRD DEGREE CORROSION|CORROS 70-79% OF BODY SURFACE W 10-19% THIRD DEGREE CORROS
C2873921|T047|E08.44|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH DIABETIC AMYOTROPHY|DIABETES DUE TO UNDERLYING CONDITION W DIABETIC AMYOTROPHY
C2882666|T047|I69.943|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING RIGHT NON-DOMINANT SIDE|MONOPLG LOW LMB FOL UNSP CEREBVASC DIS AFF RIGHT NONDOM SIDE
C2882665|T047|I69.942|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING LEFT DOMINANT SIDE|MONOPLG LOW LMB FOL UNSP CEREBVASC DISEASE AFF LEFT DOM SIDE
C2873915|T047|E08.40|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH DIABETIC NEUROPATHY, UNSPECIFIED|DIABETES DUE TO UNDERLYING CONDITION W DIABETIC NEUROP, UNSP
C2873916|T047|E08.41|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH DIABETIC MONONEUROPATHY|DIABETES DUE TO UNDRL CONDITION W DIABETIC MONONEUROPATHY
C2873918|T047|E08.42|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH DIABETIC POLYNEUROPATHY|DIABETES DUE TO UNDERLYING CONDITION W DIABETIC POLYNEUROP
C2873920|T047|E08.43|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH DIABETIC AUTONOMIC (POLY)NEUROPATHY|DIAB DUE TO UNDRL COND W DIABETIC AUTONM (POLY)NEUROPATHY
C2882668|T047|I69.949|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING UNSPECIFIED SIDE|MONOPLG LOW LMB FOL UNSP CEREBVASC DISEASE AFF UNSP SIDE
C0838545|T047|M46.83|ICD10CM|OTHER SPECIFIED INFLAMMATORY SPONDYLOPATHIES, CERVICOTHORACIC REGION|OTH INFLAMMATORY SPONDYLOPATHIES, CERVICOTHORACIC REGION
C0838551|T047|M46.80|ICD10CM|OTHER SPECIFIED INFLAMMATORY SPONDYLOPATHIES, SITE UNSPECIFIED|OTH INFLAMMATORY SPONDYLOPATHIES, SITE UNSPECIFIED
C0838543|T047|M46.81|ICD10CM|OTHER SPECIFIED INFLAMMATORY SPONDYLOPATHIES, OCCIPITO-ATLANTO-AXIAL REGION|OTH INFLAMMATORY SPONDYLOPATHIES, OCCIPT-ATLAN-AX REGION
C0838548|T047|M46.86|ICD10AM|OTHER SPECIFIED INFLAMMATORY SPONDYLOPATHIES, LUMBAR REGION|OTHER SPECIFIED INFLAMMATORY SPONDYLOPATHIES, LUMBAR REGION
C2873922|T047|E08.49|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH OTHER DIABETIC NEUROLOGICAL COMPLICATION|DIABETES DUE TO UNDRL CONDITION W OTH DIABETIC NEURO COMP
C0838546|T047|M46.84|ICD10CM|OTHER SPECIFIED INFLAMMATORY SPONDYLOPATHIES, THORACIC REGION|OTH INFLAMMATORY SPONDYLOPATHIES, THORACIC REGION
C0838547|T047|M46.85|ICD10CM|OTHER SPECIFIED INFLAMMATORY SPONDYLOPATHIES, THORACOLUMBAR REGION|OTH INFLAMMATORY SPONDYLOPATHIES, THORACOLUMBAR REGION
C2889909|T037|T82.319A|ICD10CM|BREAKDOWN (MECHANICAL) OF UNSPECIFIED VASCULAR GRAFTS, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF UNSP VASCULAR GRAFTS, INIT ENCNTR
C0494789|T047|K73.2|DMDICD10|CHRONIC ACTIVE HEPATITIS, NOT ELSEWHERE CLASSIFIED|CHRONISCHE AKTIVE HEPATITIS, ANDERENORTS NICHT KLASSIFIZIERT
C2859981|T037|S78.019S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT UNSPECIFIED HIP JOINT, SEQUELA|COMPLETE TRAUMATIC AMPUTATION AT UNSP HIP JOINT, SEQUELA
C2901299|T046|M84.564A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, LEFT FIBULA, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, LEFT FIBULA, INIT
C2887209|T047|I83.208|ICD10CM|VARICOSE VEINS OF UNSPECIFIED LOWER EXTREMITY WITH BOTH ULCER OF OTHER PART OF LOWER EXTREMITY AND INFLAMMATION|VARICOS VN UNSP LOW EXTRM W ULC OTH PRT LOW EXTRM AND INFLAM
C2887210|T047|I83.209|ICD10CM|VARICOSE VEINS OF UNSPECIFIED LOWER EXTREMITY WITH BOTH ULCER OF UNSPECIFIED SITE AND INFLAMMATION|VARICOS VN UNSP LOW EXTRM W ULC OF UNSP SITE AND INFLAM
C2859979|T037|S78.019A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT UNSPECIFIED HIP JOINT, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION AT UNSP HIP JOINT, INIT ENCNTR
C2887203|T047|I83.202|ICD10CM|VARICOSE VEINS OF UNSPECIFIED LOWER EXTREMITY WITH BOTH ULCER OF CALF AND INFLAMMATION|VARICOS VN UNSP LOW EXTRM W ULC OF CALF AND INFLAMMATION
C2887204|T047|I83.203|ICD10CM|VARICOSE VEINS OF UNSPECIFIED LOWER EXTREMITY WITH BOTH ULCER OF ANKLE AND INFLAMMATION|VARICOS VN UNSP LOW EXTRM W ULC OF ANKLE AND INFLAMMATION
C2887202|T047|I83.201|ICD10CM|VARICOSE VEINS OF UNSPECIFIED LOWER EXTREMITY WITH BOTH ULCER OF THIGH AND INFLAMMATION|VARICOS VN UNSP LOW EXTRM W ULC OF THIGH AND INFLAMMATION
C2887206|T047|I83.204|ICD10CM|VARICOSE VEINS OF UNSPECIFIED LOWER EXTREMITY WITH BOTH ULCER OF HEEL AND MIDFOOT AND INFLAMMATION|VARICOS VN UNSP LOW EXTRM W ULC OF HEEL AND MIDFT AND INFLAM
C2887208|T047|I83.205|ICD10CM|VARICOSE VEINS OF UNSPECIFIED LOWER EXTREMITY WITH BOTH ULCER OTHER PART OF FOOT AND INFLAMMATION|VARICOS VN UNSP LOW EXTRM W ULC OTH PART OF FOOT AND INFLAM
C2855984|T037|S68.519S|ICD10CM|COMPLETE TRAUMATIC TRANSPHALANGEAL AMPUTATION OF UNSPECIFIED THUMB, SEQUELA|COMPLETE TRAUMATIC TRNSPHAL AMPUTATION OF THMB, SEQUELA
C2833540|T037|S12.531B|ICD10CM|UNSPECIFIED TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP TRAUM NONDISP SPONDYLOLYSIS OF SIXTH CERVCAL VERT, 7THB
C2833539|T037|S12.531A|ICD10CM|UNSPECIFIED TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP TRAUM NONDISP SPONDYLOLYSIS OF SIXTH CERVCAL VERT, INIT
C2874404|T048|F10.29|ICD10CM|ALCOHOL DEPENDENCE WITH UNSPECIFIED ALCOHOL-INDUCED DISORDER|ALCOHOL DEPENDENCE WITH UNSPECIFIED ALCOHOL-INDUCED DISORDER
C4268209|T048|F10.26|ICD10CM|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PERSISTING AMNESTIC DISORDER|ALCOHOL USE DISORDER, SEVERE, WITH ALCOHOL-INDUCED MAJOR NEUROCOGNITIVE DISORDER, AMNESTIC-CONFABULATORY TYPE
C4268211|T048|F10.27|ICD10CM|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PERSISTING DEMENTIA|ALCOHOL USE DISORDER, SEVERE, WITH ALCOHOL-INDUCED MAJOR NEUROCOGNITIVE DISORDER, NONAMNESTIC-CONFABULATORY TYPE
C4268207|T048|F10.24|ICD10CM|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED MOOD DISORDER|ALCOHOL USE DISORDER, SEVERE, WITH ALCOHOL-INDUCED DEPRESSIVE DISORDER
C2837639|T037|S32.052A|ICD10CM|UNSTABLE BURST FRACTURE OF FIFTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSTABLE BURST FRACTURE OF FIFTH LUMBAR VERTEBRA, INIT
C4236929|T048|F10.20|ICD10CM|ALCOHOL DEPENDENCE, UNCOMPLICATED|ALCOHOL USE DISORDER, SEVERE
C4509037|T048|F10.21|ICD10CM|ALCOHOL DEPENDENCE, IN REMISSION|ALCOHOL USE DISORDER, SEVERE, IN SUSTAINED REMISSION
C2887161|T047|I82.C13|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF INTERNAL JUGULAR VEIN, BILATERAL|ACUTE EMBOLISM AND THROMBOSIS OF INT JUGULAR VEIN, BILATERAL
C2887160|T047|I82.C12|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF LEFT INTERNAL JUGULAR VEIN|ACUTE EMBOLISM AND THROMBOSIS OF LEFT INTERNAL JUGULAR VEIN
C2887159|T047|I82.C11|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF RIGHT INTERNAL JUGULAR VEIN|ACUTE EMBOLISM AND THROMBOSIS OF RIGHT INTERNAL JUGULAR VEIN
C2833465|T037|S12.430A|ICD10CM|UNSPECIFIED TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP TRAUM DISPL SPONDYLOLYSIS OF FIFTH CERVCAL VERT, INIT
C2887162|T047|I82.C19|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED INTERNAL JUGULAR VEIN|ACUTE EMBOLISM AND THROMBOSIS OF UNSP INTERNAL JUGULAR VEIN
C2901832|T047|M86.252|ICD10CM|SUBACUTE OSTEOMYELITIS, LEFT FEMUR|SUBACUTE OSTEOMYELITIS, LEFT FEMUR
C2901831|T047|M86.251|ICD10CM|SUBACUTE OSTEOMYELITIS, RIGHT FEMUR|SUBACUTE OSTEOMYELITIS, RIGHT FEMUR
C2891335|T047||ICD10CM|NECROSIS OF AMPUTATION STUMP, RIGHT UPPER EXTREMITY
C2891334|T037|T87.50|ICD10CM|NECROSIS OF AMPUTATION STUMP, UNSPECIFIED EXTREMITY|NECROSIS OF AMPUTATION STUMP, UNSPECIFIED EXTREMITY
C2891337|T047||ICD10CM|NECROSIS OF AMPUTATION STUMP, RIGHT LOWER EXTREMITY
C2901833|T047|M86.259|ICD10CM|SUBACUTE OSTEOMYELITIS, UNSPECIFIED FEMUR|SUBACUTE OSTEOMYELITIS, UNSPECIFIED FEMUR
C2886774|T037|T79.A9XA|ICD10CM|TRAUMATIC COMPARTMENT SYNDROME OF OTHER SITES, INITIAL ENCOUNTER|TRAUMATIC COMPARTMENT SYNDROME OF OTHER SITES, INIT ENCNTR
C2891338|T047||ICD10CM|NECROSIS OF AMPUTATION STUMP, LEFT LOWER EXTREMITY
C2831982|T037|S06.1X2S|ICD10CM|TRAUMATIC CEREBRAL EDEMA WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|TRAUMATIC CEREBRAL EDEMA W LOC OF 31-59 MIN, SEQUELA
C2831980|T037|S06.1X2A|ICD10CM|TRAUMATIC CEREBRAL EDEMA WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|TRAUMATIC CEREBRAL EDEMA W LOC OF 31-59 MIN, INIT
C0039236|T047|I47.9|DMDICD10|PAROXYSMAL TACHYCARDIA, UNSPECIFIED|PAROXYSMALE TACHYKARDIE, NICHT NAEHER BEZEICHNET
C0042514|T047|I47.2|DMDICD10|VENTRICULAR TACHYCARDIA|VENTRIKULAERE TACHYKARDIE
C0349069|T046|I47.0|DMDICD10|RE-ENTRY VENTRICULAR ARRHYTHMIA|VENTRIKULAERE ARRHYTHMIE DURCH RE-ENTRY
C3264368|T033|I47.1|ICD10CM|SUPRAVENTRICULAR TACHYCARDIA|ATRIOVENTRICULAR RE-ENTRANT (NODAL) TACHYCARDIA [AVNRT] [AVRT]
C2873999|T047|E09.618|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH OTHER DIABETIC ARTHROPATHY|DRUG/CHEM DIABETES MELLITUS W OTH DIABETIC ARTHROPATHY
C2874754|T048|F18.159|ICD10CM|INHALANT ABUSE WITH INHALANT-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|INHALANT ABUSE WITH INHALANT-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED
C2873998|T047|E09.610|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH DIABETIC NEUROPATHIC ARTHROPATHY|DRUG/CHEM DIABETES W DIABETIC NEUROPATHIC ARTHROPATHY
C2874753|T048|F18.151|ICD10CM|INHALANT ABUSE WITH INHALANT-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|INHALANT ABUSE W INHALNT-INDUCE PSYCH DISORDER W HALLUCIN
C2874752|T048|F18.150|ICD10CM|INHALANT ABUSE WITH INHALANT-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|INHALANT ABUSE W INHALNT-INDUCE PSYCH DISORDER W DELUSIONS
C2902438|T047|M90.542|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, LEFT HAND|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, LEFT HAND
C2833906|T037|S14.117A|ICD10CM|COMPLETE LESION AT C7 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION AT C7 LEVEL OF CERVICAL SPINAL CORD, INIT
C2859202|T037|S73.025A|ICD10CM|OBTURATOR DISLOCATION OF LEFT HIP, INITIAL ENCOUNTER|OBTURATOR DISLOCATION OF LEFT HIP, INITIAL ENCOUNTER
C2833907|T037|S14.117D|ICD10CM|COMPLETE LESION AT C7 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION AT C7 LEVEL OF CERVICAL SPINAL CORD, SUBS
C2910347|T047|Q87.42|ICD10CM|MARFAN'S SYNDROME WITH OCULAR MANIFESTATIONS|MARFAN'S SYNDROME WITH OCULAR MANIFESTATIONS
C0039445|T047|I78.0|DMDICD10|HEREDITARY HEMORRHAGIC TELANGIECTASIA|HEREDITAERE HAEMORRHAGISCHE TELEANGIEKTASIE
C2890674|T037|T84.194A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTERNAL FIXATION DEVICE OF RIGHT FEMUR, INITIAL ENCOUNTER|MECH COMPL OF INTERNAL FIXATION DEVICE OF RIGHT FEMUR, INIT
C2889583|T047|M08.43|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED WRIST|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, WRIST
C2856107|T037|S68.729A|ICD10CM|PARTIAL TRAUMATIC TRANSMETACARPAL AMPUTATION OF UNSPECIFIED HAND, INITIAL ENCOUNTER|PARTIAL TRAUMATIC TRANSMETCRPL AMPUTATION OF UNSP HAND, INIT
C2889581|T047|M08.431|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, RIGHT WRIST|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, RIGHT WRIST
C2889582|T047|M08.432|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, LEFT WRIST|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, LEFT WRIST
C0348694|T047|J62.8|DMDICD10|PNEUMOCONIOSIS DUE TO OTHER DUST CONTAINING SILICA|PNEUMOKONIOSE DURCH SONSTIGEN QUARZSTAUB
C2856846|T037|S72.044C|ICD10CM|NONDISPLACED FRACTURE OF BASE OF NECK OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF BASE OF NK OF R FEMR, 7THC
C2856845|T037|S72.044B|ICD10CM|NONDISPLACED FRACTURE OF BASE OF NECK OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF BASE OF NK OF R FEMR, INIT FOR OPN FX TYPE I/2
C2856844|T037|S72.044A|ICD10CM|NONDISPLACED FRACTURE OF BASE OF NECK OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF BASE OF NECK OF RIGHT FEMUR, INIT FOR CLOS FX
C2832588|T037|S06.819S|ICD10CM|INJURY OF RIGHT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|INJ R INT CAROTID, INTCR W LOC OF UNSP DURATION, SEQUELA
C0238377|T047|J62.0|DMDICD10|PNEUMOCONIOSIS DUE TO TALC DUST|PNEUMOKONIOSE DURCH TALKUM-STAUB
C2843342|T037|S48.929A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED SHOULDER AND UPPER ARM, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP OF UNSP SHLDR/UP ARM, LEVEL UNSP, INIT
C2857961|T037|S72.343C|ICD10CM|DISPLACED SPIRAL FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL SPIRAL FX SHAFT OF UNSP FEMR, 7THC
C2857960|T037|S72.343B|ICD10CM|DISPLACED SPIRAL FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL SPIRAL FX SHAFT OF UNSP FEMR, INIT FOR OPN FX TYPE I/2
C2857959|T037|S72.343A|ICD10CM|DISPLACED SPIRAL FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED SPIRAL FRACTURE OF SHAFT OF UNSP FEMUR, INIT
C2833346|T037|S12.24XB|ICD10CM|TYPE III TRAUMATIC SPONDYLOLISTHESIS OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE III TRAUM SPONDYLOLYSIS OF 3RD CERVCAL VERT, 7THB
C2833345|T037|S12.24XA|ICD10CM|TYPE III TRAUMATIC SPONDYLOLISTHESIS OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE III TRAUM SPONDYLOLYSIS OF THIRD CERVCAL VERTEBRA, INIT
C2889158|T047|M05.169|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP KNEE
C4268213|T048|F10.288|ICD10CM|ALCOHOL DEPENDENCE WITH OTHER ALCOHOL-INDUCED DISORDER|ALCOHOL USE DISORDER, SEVERE, WITH ALCOHOL-INDUCED MILD NEUROCOGNITIVE DISORDER
C2889156|T047|M05.161|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT KNEE|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2858491|T037|S72.424A|ICD10CM|NONDISPLACED FRACTURE OF LATERAL CONDYLE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF LATERAL CONDYLE OF RIGHT FEMUR, INIT
C2889157|T047|M05.162|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT KNEE|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT KNEE
C2874402|T048|F10.282|ICD10CM|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED SLEEP DISORDER|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED SLEEP DISORDER
C2874401|T048|F10.281|ICD10CM|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED SEXUAL DYSFUNCTION|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED SEXUAL DYSFUNCTION
C2874400|T048|F10.280|ICD10CM|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED ANXIETY DISORDER|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED ANXIETY DISORDER
C2901835|T047|M86.262|ICD10CM|SUBACUTE OSTEOMYELITIS, LEFT TIBIA AND FIBULA|SUBACUTE OSTEOMYELITIS, LEFT TIBIA AND FIBULA
C2835363|T037|S22.059B|ICD10CM|UNSPECIFIED FRACTURE OF T5-T6 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF T5-T6 VERTEBRA, INIT FOR OPN FX
C2901834|T047|M86.261|ICD10CM|SUBACUTE OSTEOMYELITIS, RIGHT TIBIA AND FIBULA|SUBACUTE OSTEOMYELITIS, RIGHT TIBIA AND FIBULA
C2835362|T037|S22.059A|ICD10CM|UNSPECIFIED FRACTURE OF T5-T6 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF T5-T6 VERTEBRA, INIT FOR CLOS FX
C4268627|T047|K55.049|ICD10CM|ACUTE INFARCTION OF LARGE INTESTINE, EXTENT UNSPECIFIED|ACUTE INFARCTION OF LARGE INTESTINE, EXTENT UNSPECIFIED
C4268625|T047|K55.041|ICD10CM|FOCAL (SEGMENTAL) ACUTE INFARCTION OF LARGE INTESTINE|FOCAL (SEGMENTAL) ACUTE INFARCTION OF LARGE INTESTINE
C4268626|T047||ICD10CM|DIFFUSE ACUTE INFARCTION OF LARGE INTESTINE
C2835798|T037|S24.131D|ICD10CM|ANTERIOR CORD SYNDROME AT T1 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|ANTERIOR CORD SYNDROME AT T1, SUBS
C2530958|T061|D704|ICD10PCS|CYCLIC NEUTROPENIA|RADIATION THERAPY @ LYMPHATIC AND HEMATOLOGIC SYSTEM @ BEAM RADIATION @ LYMPHATICS, AXILLARY
C2530945|T061|D703|ICD10PCS|NEUTROPENIA DUE TO INFECTION|RADIATION THERAPY @ LYMPHATIC AND HEMATOLOGIC SYSTEM @ BEAM RADIATION @ LYMPHATICS, NECK
C2873811|T046|D70.2|ICD10CM|OTHER DRUG-INDUCED AGRANULOCYTOSIS|OTHER DRUG-INDUCED AGRANULOCYTOSIS
C2883114|T046|I82.492|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF OTHER SPECIFIED DEEP VEIN OF LEFT LOWER EXTREMITY|ACUTE EMBOLISM AND THROMBOSIS OF DEEP VEIN OF L LOW EXTREM
C2883115|T046|I82.493|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF OTHER SPECIFIED DEEP VEIN OF LOWER EXTREMITY, BILATERAL|ACUTE EMBOLISM AND THOMBOS OF DEEP VEIN OF LOW EXTRM, BI
C2874943|T033|F40.233|ICD10CM|FEAR OF INJURY|FEAR OF INJURY
C2874942|T048|F40.232|ICD10CM|FEAR OF OTHER MEDICAL CARE|FEAR OF OTHER MEDICAL CARE
C2874941|T048|F40.231|ICD10CM|FEAR OF INJECTIONS AND TRANSFUSIONS|FEAR OF INJECTIONS AND TRANSFUSIONS
C0522183|T048|F40.230|ICD10CM|FEAR OF BLOOD|FEAR OF BLOOD
C2883116|T046|I82.499|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF OTHER SPECIFIED DEEP VEIN OF UNSPECIFIED LOWER EXTREMITY|ACUTE EMBOLISM AND THROMBOSIS OF DEEP VEIN OF UNSP LOW EXTRM
C0027947|T047|D70.9|ICD10CM|NEUTROPENIA, UNSPECIFIED|NEUTROPENIA, UNSPECIFIED
C3263991|T047|G40.A01|ICD10CM|ABSENCE EPILEPTIC SYNDROME, NOT INTRACTABLE, WITH STATUS EPILEPTICUS|ABSENCE EPILEPTIC SYNDROME, NOT INTRACTABLE, W STAT EPI
C2884086|T037|T52.0X2A|ICD10CM|TOXIC EFFECT OF PETROLEUM PRODUCTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF PETROLEUM PRODUCTS, SELF-HARM, INIT
C4269508|T037|S02.640S|ICD10CM|FRACTURE OF RAMUS OF MANDIBLE, UNSPECIFIED SIDE, SEQUELA|FRACTURE OF RAMUS OF MANDIBLE, UNSPECIFIED SIDE, SEQUELA
C0751394|T191||ICD10CM|MALIGNANT NEOPLASM OF HEAD, FACE AND NECK
C1998032|T191||ICD10CM|MALIGNANT NEOPLASM OF THORAX
C0153662|T191|C76.2|DMDICD10|MALIGNANT NEOPLASM OF ABDOMEN|BOESARTIGE NEUBILDUNG UNGENAU BEZEICHNETER LOKALISATIONEN: ABDOMEN
C3665513|T191||ICD10CM|MALIGNANT NEOPLASM OF PELVIS
C2858765|T037|S72.452A|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPL SUPRCNDL FX W/O INTRCNDL EXTN LOWER END L FEMUR, INIT
C2858766|T037|S72.452B|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL SUPRCNDL FX W/O INTRCNDL EXTN LOW END L FEMR, 7THB
C2858767|T037|S72.452C|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL SUPRCNDL FX W/O INTRCNDL EXTN LOW END L FEMR, 7THC
C2977945|T191|C76.8|ICD10CM|MALIGNANT NEOPLASM OF OTHER SPECIFIED ILL-DEFINED SITES|MALIGNANT NEOPLASM OF OTHER SPECIFIED ILL-DEFINED SITES
C2875183|T047|G43.819|ICD10CM|OTHER MIGRAINE, INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|OTHER MIGRAINE, INTRACTABLE, WITHOUT STATUS MIGRAINOSUS
C2884088|T037|T52.0X2S|ICD10CM|TOXIC EFFECT OF PETROLEUM PRODUCTS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF PETROLEUM PRODUCTS, SELF-HARM, SEQUELA
C2832093|T037|S06.309S|ICD10CM|UNSPECIFIED FOCAL TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|UNSP FOCAL TBI W LOC OF UNSP DURATION, SEQUELA
C0837507|T047|M05.09|ICD10CM|FELTY'S SYNDROME, MULTIPLE SITES|FELTY'S SYNDROME, MULTIPLE SITES
C2832091|T037|S06.309A|ICD10CM|UNSPECIFIED FOCAL TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|UNSP FOCAL TBI W LOC OF UNSP DURATION, INIT
C4268062|T047|E10.3599|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|TYPE 1 DIAB WITH PROLIF DIAB RTNOP WITHOUT MCLR EDEMA, UNSP
C2883045|T047|I75.019|ICD10CM|ATHEROEMBOLISM OF UNSPECIFIED UPPER EXTREMITY|ATHEROEMBOLISM OF UNSPECIFIED UPPER EXTREMITY
C4268060|T047|E10.3592|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|TYPE 1 DIAB WITH PROLIF DIAB RTNOP WITHOUT MCLR EDEMA, L EYE
C4268061|T047|E10.3593|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|TYPE 1 DIAB WITH PROLIF DIAB RTNOP WITHOUT MACULAR EDEMA, BI
C4268059|T047|E10.3591|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|TYPE 1 DIAB WITH PROLIF DIAB RTNOP WITHOUT MCLR EDEMA, R EYE
C2883043|T047|I75.012|ICD10CM|ATHEROEMBOLISM OF LEFT UPPER EXTREMITY|ATHEROEMBOLISM OF LEFT UPPER EXTREMITY
C2883044|T047|I75.013|ICD10CM|ATHEROEMBOLISM OF BILATERAL UPPER EXTREMITIES|ATHEROEMBOLISM OF BILATERAL UPPER EXTREMITIES
C2883042|T047|I75.011|ICD10CM|ATHEROEMBOLISM OF RIGHT UPPER EXTREMITY|ATHEROEMBOLISM OF RIGHT UPPER EXTREMITY
C2890596|T037|T84.114A|ICD10CM|BREAKDOWN (MECHANICAL) OF INTERNAL FIXATION DEVICE OF RIGHT FEMUR, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF INT FIX OF RIGHT FEMUR, INIT
C2860040|T037|S78.922A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT HIP AND THIGH, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|PARTIAL TRAUM AMP OF LEFT HIP AND THIGH, LEVEL UNSP, INIT
C2900932|T046|M84.434A|ICD10CM|PATHOLOGICAL FRACTURE, LEFT RADIUS, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, LEFT RADIUS, INIT ENCNTR FOR FRACTURE
C2860041|T037|S78.922D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT HIP AND THIGH, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|PARTIAL TRAUM AMP OF LEFT HIP AND THIGH, LEVEL UNSP, SUBS
C2889067|T047|M02.352|ICD10CM|REITER'S DISEASE, LEFT HIP|REITER'S DISEASE, LEFT HIP
C2889066|T047|M02.351|ICD10CM|REITER'S DISEASE, RIGHT HIP|REITER'S DISEASE, RIGHT HIP
C2860042|T037|S78.922S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT HIP AND THIGH, LEVEL UNSPECIFIED, SEQUELA|PARTIAL TRAUM AMP OF LEFT HIP AND THIGH, LEVEL UNSP, SEQUELA
C2889068|T047|M02.359|ICD10CM|REITER'S DISEASE, UNSPECIFIED HIP|REITER'S DISEASE, UNSPECIFIED HIP
C2884448|T037|T55.1X2S|ICD10CM|TOXIC EFFECT OF DETERGENTS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF DETERGENTS, INTENTIONAL SELF-HARM, SEQUELA
C2977870|T037|S32.592B|ICD10CM|OTHER SPECIFIED FRACTURE OF LEFT PUBIS, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF LEFT PUBIS, INIT ENCNTR FOR OPEN FRACTURE
C3264040|T047|G43.B1|ICD10CM|OPHTHALMOPLEGIC MIGRAINE, INTRACTABLE|OPHTHALMOPLEGIC MIGRAINE, WITH REFRACTORY MIGRAINE
C3264039|T047|G43.B0|ICD10CM|OPHTHALMOPLEGIC MIGRAINE, NOT INTRACTABLE|OPHTHALMOPLEGIC MIGRAINE, WITHOUT REFRACTORY MIGRAINE
C2843275|T037|S48.012S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEFT SHOULDER JOINT, SEQUELA|COMPLETE TRAUMATIC AMPUTATION AT L SHOULDER JT, SEQUELA
C2832204|T037|S06.336S|ICD10CM|CONTUSION AND LACERATION OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|CONTUS/LAC CEREB, W LOC >24 HR W/O RET CONSC W SURV, SEQUELA
C2901973|T046|M87.066|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED FIBULA|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED FIBULA
C2835190|T037|S22.010A|ICD10CM|WEDGE COMPRESSION FRACTURE OF FIRST THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|WEDGE COMPRESSION FRACTURE OF FIRST THORACIC VERTEBRA, INIT
C2835191|T037|S22.010B|ICD10CM|WEDGE COMPRESSION FRACTURE OF FIRST THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|WEDGE COMPRSN FX FIRST THOR VERTEBRA, INIT FOR OPN FX
C2843273|T037|S48.012A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEFT SHOULDER JOINT, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION AT LEFT SHOULDER JOINT, INIT
C2832202|T037|S06.336A|ICD10CM|CONTUSION AND LACERATION OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|CONTUS/LAC CEREB, W LOC >24 HR W/O RET CONSC W SURV, INIT
C0153434|T191|C18.4|DMDICD10|MALIGNANT NEOPLASM OF TRANSVERSE COLON|BOESARTIGE NEUBILDUNG: COLON TRANSVERSUM
C0153440|T191|C18.5|DMDICD10|MALIGNANT NEOPLASM OF SPLENIC FLEXURE|BOESARTIGE NEUBILDUNG: FLEXURA COLI SINISTRA [LIENALIS]
C0153435|T191|C18.6|DMDICD10|MALIGNANT NEOPLASM OF DESCENDING COLON|BOESARTIGE NEUBILDUNG: COLON DESCENDENS
C0864870|T191|C18.7|ICD10CM|MALIGNANT NEOPLASM OF SIGMOID COLON|MALIGNANT NEOPLASM OF SIGMOID (FLEXURE)
C2874462|T048|F11.950|ICD10CM|OPIOID USE, UNSPECIFIED WITH OPIOID-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|OPIOID USE, UNSP W OPIOID-INDUC PSYCH DISORDER W DELUSIONS
C0496779|T191|C18.1|DMDICD10|MALIGNANT NEOPLASM OF APPENDIX|BOESARTIGE NEUBILDUNG: APPENDIX VERMIFORMIS
C0348384|T191|C78.8|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF OTHER DIGESTIVE ORGANS|SECONDARY MALIGNANT NEOPLASM OF OTHER AND UNSPECIFIED DIGESTIVE ORGANS
C0153433|T191|C18.3|DMDICD10|MALIGNANT NEOPLASM OF HEPATIC FLEXURE|BOESARTIGE NEUBILDUNG: FLEXURA COLI DEXTRA [HEPATICA]
C0349051|T191|C18.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF COLON|BOESARTIGE NEUBILDUNG: KOLON, MEHRERE TEILBEREICHE UEBERLAPPEND
C2874464|T048|F11.959|ICD10CM|OPIOID USE, UNSPECIFIED WITH OPIOID-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|OPIOID USE, UNSP W OPIOID-INDUCED PSYCHOTIC DISORDER, UNSP
C2845962|T191|C78.80|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF UNSPECIFIED DIGESTIVE ORGAN|SECONDARY MALIGNANT NEOPLASM OF UNSPECIFIED DIGESTIVE ORGAN
C2886921|T037|T81.512S|ICD10CM|ADHESIONS DUE TO FOREIGN BODY ACCIDENTALLY LEFT IN BODY FOLLOWING KIDNEY DIALYSIS, SEQUELA|ADHES DUE TO FB ACC LEFT IN BODY FOL KIDNEY DIALYSIS, SQLA
C2905652|T037|X71.1XXS|ICD10CM|INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION WHILE IN SWIMMING POOL, SEQUELA|SELF-HARM BY DROWN WHILE IN SWIMMING POOL, SEQUELA
C2883787|T037|T50.992S|ICD10CM|POISONING BY OTHER DRUGS, MEDICAMENTS AND BIOLOGICAL SUBSTANCES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH DRUG/MEDS/BIOL SUBST, SELF-HARM, SEQUELA
C2874221|T047|E46|ICD10CM|UNSPECIFIED PROTEIN-CALORIE MALNUTRITION|PROTEIN-CALORIE IMBALANCE NOS
C2874654|T048|F15.251|ICD10CM|OTHER STIMULANT DEPENDENCE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|OTH STIMULANT DEPEND W STIM-INDUCE PSYCH DISORDER W HALLUCIN
C2874653|T048|F15.250|ICD10CM|OTHER STIMULANT DEPENDENCE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|OTH STIM DEPEND W STIM-INDUCE PSYCH DISORDER W DELUSIONS
C2874655|T048|F15.25|ICD10CM|OTHER STIMULANT DEPENDENCE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|OTHER STIMULANT DEPENDENCE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER
C2884446|T037|T55.1X2A|ICD10CM|TOXIC EFFECT OF DETERGENTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF DETERGENTS, INTENTIONAL SELF-HARM, INIT
C2884964|T037|T59.812S|ICD10CM|TOXIC EFFECT OF SMOKE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF SMOKE, INTENTIONAL SELF-HARM, SEQUELA
C4270338|T046|T83.592A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INDWELLING URETERAL STENT, INITIAL ENCOUNTER|I/I REACT D/T INDWELLING URETERAL STENT, INITIAL ENCOUNTER
C2886961|T037|T81.522D|ICD10CM|OBSTRUCTION DUE TO FOREIGN BODY ACCIDENTALLY LEFT IN BODY FOLLOWING KIDNEY DIALYSIS, SUBSEQUENT ENCOUNTER|OBST DUE TO FB ACC LEFT IN BODY FOL KIDNEY DIALYSIS, SUBS
C2843290|T037|S48.029A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT UNSPECIFIED SHOULDER JOINT, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION AT UNSP SHOULDER JOINT, INIT
C2884336|T037|T53.92XS|ICD10CM|TOXIC EFFECT OF UNSPECIFIED HALOGEN DERIVATIVES OF ALIPHATIC AND AROMATIC HYDROCARBONS, INTENTIONAL SELF-HARM, SEQUELA|TOX EFF OF UNSP HALGN DERIV OF AROMAT HYDROCRB,SLF-HRM, SQLA
C2895193|T047|M33.92|ICD10CM|DERMATOPOLYMYOSITIS, UNSPECIFIED WITH MYOPATHY|DERMATOPOLYMYOSITIS, UNSPECIFIED WITH MYOPATHY
C2875093|T047|G40.209|ICD10CM|LOCALIZATION-RELATED (FOCAL) (PARTIAL) SYMPTOMATIC EPILEPSY AND EPILEPTIC SYNDROMES WITH COMPLEX PARTIAL SEIZURES, NOT INTRACTABLE, WITHOUT STATUS EPILEPTICUS|LOCAL-REL SYMPTC EPI W CMPLX PRT SEIZ,NOT NTRCT,W/O STAT EPI
C2838186|T037|S32.452A|ICD10CM|DISPLACED TRANSVERSE FRACTURE OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED TRANSVERSE FRACTURE OF LEFT ACETABULUM, INIT
C2838187|T037|S32.452B|ICD10CM|DISPLACED TRANSVERSE FRACTURE OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISPLACED TRANSVERSE FX LEFT ACETABULUM, INIT FOR OPN FX
C2886960|T037|T81.522A|ICD10CM|OBSTRUCTION DUE TO FOREIGN BODY ACCIDENTALLY LEFT IN BODY FOLLOWING KIDNEY DIALYSIS, INITIAL ENCOUNTER|OBST DUE TO FB ACC LEFT IN BODY FOL KIDNEY DIALYSIS, INIT
C2905651|T037|X71.1XXD|ICD10CM|INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION WHILE IN SWIMMING POOL, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY DROWN WHILE IN SWIMMING POOL, SUBS
C2877997|T037|T41.42XS|ICD10CM|POISONING BY UNSPECIFIED ANESTHETIC, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY UNSP ANESTHETIC, INTENTIONAL SELF-HARM, SEQUELA
C2884897|T037|T59.4X2A|ICD10CM|TOXIC EFFECT OF CHLORINE GAS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CHLORINE GAS, INTENTIONAL SELF-HARM, INIT
C0042510|T047||ICD10CM|VENTRICULAR FIBRILLATION
C0152173|T047||ICD10CM|VENTRICULAR FLUTTER
C2835407|T037|S22.070B|ICD10CM|WEDGE COMPRESSION FRACTURE OF T9-T10 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|WEDGE COMPRSN FRACTURE OF T9-T10 VERTEBRA, INIT FOR OPN FX
C2884899|T037|T59.4X2S|ICD10CM|TOXIC EFFECT OF CHLORINE GAS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CHLORINE GAS, INTENTIONAL SELF-HARM, SEQUELA
C2886412|T037|T71.162A|ICD10CM|ASPHYXIATION DUE TO HANGING, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|ASPHYXIATION DUE TO HANGING, INTENTIONAL SELF-HARM, INIT
C2889946|T037|T82.338A|ICD10CM|LEAKAGE OF OTHER VASCULAR GRAFTS, INITIAL ENCOUNTER|LEAKAGE OF OTHER VASCULAR GRAFTS, INITIAL ENCOUNTER
C4268167|T047|E13.3549|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, UNSPECIFIED EYE|OTH DIAB WITH PROLIF DIABETIC RTNOP WITH COMB DETACH, UNSP
C4268165|T047|E13.3542|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, LEFT EYE|OTH DIAB WITH PROLIF DIAB RTNOP WITH COMB DETACH, LEFT EYE
C4268166|T047|E13.3543|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, BILATERAL|OTH DIABETES WITH PROLIF DIABETIC RTNOP WITH COMB DETACH, BI
C4268164|T047|E13.3541|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, RIGHT EYE|OTH DIAB WITH PROLIF DIABETIC RTNOP WITH COMB DETACH, R EYE
C2835406|T037|S22.070A|ICD10CM|WEDGE COMPRESSION FRACTURE OF T9-T10 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|WEDGE COMPRESSION FRACTURE OF T9-T10 VERTEBRA, INIT
C2886414|T037|T71.162S|ICD10CM|ASPHYXIATION DUE TO HANGING, INTENTIONAL SELF-HARM, SEQUELA|ASPHYXIATION DUE TO HANGING, INTENTIONAL SELF-HARM, SEQUELA
C2911576|T033|Z99.12|ICD10CM|ENCOUNTER FOR RESPIRATOR [VENTILATOR] DEPENDENCE DURING POWER FAILURE|ENCOUNTER FOR RESPIRATOR DEPENDENCE DURING POWER FAILURE
C2911575|T033|Z99.11|ICD10CM|DEPENDENCE ON RESPIRATOR [VENTILATOR] STATUS|DEPENDENCE ON RESPIRATOR [VENTILATOR] STATUS
C2838352|T037|S32.491B|ICD10CM|OTHER SPECIFIED FRACTURE OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF RIGHT ACETABULUM, INIT FOR OPN FX
C2882886|T047|I70.538|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF OTHER PART OF LOWER LEG|ATHSCL NONAUT BIO BYPASS OF R LEG W ULCER OTH PRT LOW LEG
C2882887|T047|I70.539|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF UNSPECIFIED SITE|ATHSCL NONAUT BIO BYPASS OF RIGHT LEG W ULCER OF UNSP SITE
C2888476|T047|L89.44|ICD10CM|PRESSURE ULCER OF CONTIGUOUS SITE OF BACK, BUTTOCK AND HIP, STAGE 4|PRESSR ULCER OF CONTIG SITE OF BACK, BUTTOCK AND HIP, STG 4
C2888477|T047|L89.45|ICD10CM|PRESSURE ULCER OF CONTIGUOUS SITE OF BACK, BUTTOCK AND HIP, UNSTAGEABLE|PRESSR ULC OF CONTIG SITE OF BACK,BUTTOCK & HIP, UNSTAGEABLE
C2882883|T047|I70.534|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF HEEL AND MIDFOOT|ATHSCL NONAUT BIO BYPASS OF R LEG W ULCER OF HEEL AND MIDFT
C2882885|T047|I70.535|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF OTHER PART OF FOOT|ATHSCL NONAUT BIO BYPASS OF RIGHT LEG W ULCER OTH PRT FOOT
C2888464|T047|L89.40|ICD10CM|PRESSURE ULCER OF CONTIGUOUS SITE OF BACK, BUTTOCK AND HIP, UNSPECIFIED STAGE|PRESSR ULC OF CONTIG SITE OF BACK, BUTTOCK AND HIP, UNSP STG
C2888467|T047|L89.41|ICD10CM|PRESSURE ULCER OF CONTIGUOUS SITE OF BACK, BUTTOCK AND HIP, STAGE 1|PRESSR ULCER OF CONTIG SITE OF BACK, BUTTOCK AND HIP, STG 1
C2888470|T047|L89.42|ICD10CM|PRESSURE ULCER OF CONTIGUOUS SITE OF BACK, BUTTOCK AND HIP, STAGE 2|PRESSR ULCER OF CONTIG SITE OF BACK, BUTTOCK AND HIP, STG 2
C2888473|T047|L89.43|ICD10CM|PRESSURE ULCER OF CONTIGUOUS SITE OF BACK, BUTTOCK AND HIP, STAGE 3|PRESSR ULCER OF CONTIG SITE OF BACK, BUTTOCK AND HIP, STG 3
C2893652|T047|M12.072|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], LEFT ANKLE AND FOOT|CHRONIC POSTRHEUMATIC ARTHROPATHY, LEFT ANKLE AND FOOT
C2893651|T047|M12.071|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], RIGHT ANKLE AND FOOT|CHRONIC POSTRHEUMATIC ARTHROPATHY, RIGHT ANKLE AND FOOT
C2853954|T191|C83.98|ICD10CM|NON-FOLLICULAR (DIFFUSE) LYMPHOMA, UNSPECIFIED, LYMPH NODES OF MULTIPLE SITES|NON-FOLLIC (DIFFUSE) LYMPHOMA, UNSP, LYMPH NODES MULT SITE
C2853955|T191|C83.99|ICD10CM|NON-FOLLICULAR (DIFFUSE) LYMPHOMA, UNSPECIFIED, EXTRANODAL AND SOLID ORGAN SITES|NON-FOLLIC LYMPHOMA, UNSP, EXTRNOD AND SOLID ORGAN SITES
C2853952|T191|C83.96|ICD10CM|NON-FOLLICULAR (DIFFUSE) LYMPHOMA, UNSPECIFIED, INTRAPELVIC LYMPH NODES|NON-FOLLIC (DIFFUSE) LYMPHOMA, UNSP, INTRAPELVIC LYMPH NODES
C2853953|T191|C83.97|ICD10CM|NON-FOLLICULAR (DIFFUSE) LYMPHOMA, UNSPECIFIED, SPLEEN|NON-FOLLICULAR (DIFFUSE) LYMPHOMA, UNSPECIFIED, SPLEEN
C2853950|T191|C83.94|ICD10CM|NON-FOLLICULAR (DIFFUSE) LYMPHOMA, UNSPECIFIED, LYMPH NODES OF AXILLA AND UPPER LIMB|NON-FOLLIC LYMPHOMA, UNSP, NODES OF AXILLA AND UPPER LIMB
C2853951|T191|C83.95|ICD10CM|NON-FOLLICULAR (DIFFUSE) LYMPHOMA, UNSPECIFIED, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|NON-FOLLIC LYMPH, UNSP, NODES OF ING REGION AND LOWER LIMB
C2853948|T191|C83.92|ICD10CM|NON-FOLLICULAR (DIFFUSE) LYMPHOMA, UNSPECIFIED, INTRATHORACIC LYMPH NODES|NON-FOLLIC (DIFFUSE) LYMPHOMA, UNSP, INTRATHORAC LYMPH NODES
C2853949|T191|C83.93|ICD10CM|NON-FOLLICULAR (DIFFUSE) LYMPHOMA, UNSPECIFIED, INTRA-ABDOMINAL LYMPH NODES|NON-FOLLIC (DIFFUSE) LYMPHOMA, UNSP, INTRA-ABD LYMPH NODES
C2853946|T191|C83.90|ICD10CM|NON-FOLLICULAR (DIFFUSE) LYMPHOMA, UNSPECIFIED, UNSPECIFIED SITE|NON-FOLLICULAR (DIFFUSE) LYMPHOMA, UNSP, UNSPECIFIED SITE
C2853947|T191|C83.91|ICD10CM|NON-FOLLICULAR (DIFFUSE) LYMPHOMA, UNSPECIFIED, LYMPH NODES OF HEAD, FACE, AND NECK|NON-FOLLIC LYMPHOMA, UNSP, NODES OF HEAD, FACE, AND NECK
C2896742|T046|M80.849A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, UNSPECIFIED HAND, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, UNSP HAND, INIT
C4269424|T037|S02.600S|ICD10CM|FRACTURE OF UNSPECIFIED PART OF BODY OF MANDIBLE, UNSPECIFIED SIDE, SEQUELA|FX UNSP PART OF BODY OF MANDIBLE, UNSPECIFIED SIDE, SEQUELA
C2876201|T037|T32.55|ICD10CM|CORROSIONS INVOLVING 50-59% OF BODY SURFACE WITH 50-59% THIRD DEGREE CORROSION|CORROS 50-59% OF BODY SURFACE W 50-59% THIRD DEGREE CORROS
C2876200|T037|T32.54|ICD10CM|CORROSIONS INVOLVING 50-59% OF BODY SURFACE WITH 40-49% THIRD DEGREE CORROSION|CORROS 50-59% OF BODY SURFACE W 40-49% THIRD DEGREE CORROS
C2876197|T037|T32.51|ICD10CM|CORROSIONS INVOLVING 50-59% OF BODY SURFACE WITH 10-19% THIRD DEGREE CORROSION|CORROS 50-59% OF BODY SURFACE W 10-19% THIRD DEGREE CORROS
C2876199|T037|T32.53|ICD10CM|CORROSIONS INVOLVING 50-59% OF BODY SURFACE WITH 30-39% THIRD DEGREE CORROSION|CORROS 50-59% OF BODY SURFACE W 30-39% THIRD DEGREE CORROS
C2876198|T037|T32.52|ICD10CM|CORROSIONS INVOLVING 50-59% OF BODY SURFACE WITH 20-29% THIRD DEGREE CORROSION|CORROS 50-59% OF BODY SURFACE W 20-29% THIRD DEGREE CORROS
C2869887|T037|S98.911A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT FOOT, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMP OF RIGHT FOOT, LEVEL UNSP, INIT
C2885027|T037|T60.1X2A|ICD10CM|TOXIC EFFECT OF HALOGENATED INSECTICIDES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF HALOGENATED INSECTICIDES, SELF-HARM, INIT
C1701940|T047||ICD10CM|VENTILATOR ASSOCIATED PNEUMONIA
C2228900|T046|J95.850|ICD10CM|MECHANICAL COMPLICATION OF RESPIRATOR|MECHANICAL COMPLICATION OF RESPIRATOR
C2905713|T037|X74.8XXD|ICD10CM|INTENTIONAL SELF-HARM BY OTHER FIREARM DISCHARGE, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY OTH FIREARM DISCHARGE, SUBS ENCNTR
C2905712|T037|X74.8XXA|ICD10CM|INTENTIONAL SELF-HARM BY OTHER FIREARM DISCHARGE, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY OTH FIREARM DISCHARGE, INIT ENCNTR
C2887509|T047|J95.859|ICD10CM|OTHER COMPLICATION OF RESPIRATOR [VENTILATOR]|OTHER COMPLICATION OF RESPIRATOR [VENTILATOR]
C2905658|T037|X71.3XXA|ICD10CM|INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION IN NATURAL WATER, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY DROWN IN NATURAL WATER, INIT
C2905659|T037|X71.3XXD|ICD10CM|INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION IN NATURAL WATER, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY DROWN IN NATURAL WATER, SUBS
C2854021|T191|C84.Z8|ICD10CM|OTHER MATURE T/NK-CELL LYMPHOMAS, LYMPH NODES OF MULTIPLE SITES|OTH MATURE T/NK-CELL LYMPHOMAS, LYMPH NODES MULT SITE
C2854022|T191|C84.Z9|ICD10CM|OTHER MATURE T/NK-CELL LYMPHOMAS, EXTRANODAL AND SOLID ORGAN SITES|OTH MATURE T/NK-CELL LYMPH, EXTRNOD AND SOLID ORGAN SITES
C2905714|T037|X74.8XXS|ICD10CM|INTENTIONAL SELF-HARM BY OTHER FIREARM DISCHARGE, SEQUELA|INTENTIONAL SELF-HARM BY OTHER FIREARM DISCHARGE, SEQUELA
C2874623|T048|F14.99|ICD10CM|COCAINE USE, UNSPECIFIED WITH UNSPECIFIED COCAINE-INDUCED DISORDER|COCAINE USE, UNSP WITH UNSPECIFIED COCAINE-INDUCED DISORDER
C2854013|T191|C84.Z0|ICD10CM|OTHER MATURE T/NK-CELL LYMPHOMAS, UNSPECIFIED SITE|OTHER MATURE T/NK-CELL LYMPHOMAS, UNSPECIFIED SITE
C2854014|T191|C84.Z1|ICD10CM|OTHER MATURE T/NK-CELL LYMPHOMAS, LYMPH NODES OF HEAD, FACE, AND NECK|OTH MATURE T/NK-CELL LYMPH, NODES OF HEAD, FACE, AND NECK
C2854015|T191|C84.Z2|ICD10CM|OTHER MATURE T/NK-CELL LYMPHOMAS, INTRATHORACIC LYMPH NODES|OTHER MATURE T/NK-CELL LYMPHOMAS, INTRATHORACIC LYMPH NODES
C2854016|T191|C84.Z3|ICD10CM|OTHER MATURE T/NK-CELL LYMPHOMAS, INTRA-ABDOMINAL LYMPH NODES|OTH MATURE T/NK-CELL LYMPHOMAS, INTRA-ABDOMINAL LYMPH NODES
C2854017|T191|C84.Z4|ICD10CM|OTHER MATURE T/NK-CELL LYMPHOMAS, LYMPH NODES OF AXILLA AND UPPER LIMB|OTH MATURE T/NK-CELL LYMPH, NODES OF AXILLA AND UPPER LIMB
C2854018|T191|C84.Z5|ICD10CM|OTHER MATURE T/NK-CELL LYMPHOMAS, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|OTH MATURE T/NK-CELL LYMPH, NODES OF ING RGN AND LOWER LIMB
C2854019|T191|C84.Z6|ICD10CM|OTHER MATURE T/NK-CELL LYMPHOMAS, INTRAPELVIC LYMPH NODES|OTHER MATURE T/NK-CELL LYMPHOMAS, INTRAPELVIC LYMPH NODES
C2854020|T191|C84.Z7|ICD10CM|OTHER MATURE T/NK-CELL LYMPHOMAS, SPLEEN|OTHER MATURE T/NK-CELL LYMPHOMAS, SPLEEN
C0349208|T048|F30|DMDICD10|MANIC EPISODE, UNSPECIFIED|MANISCHE EPISODE
C0349207|T048|F30.8|DMDICD10|OTHER MANIC EPISODES|SONSTIGE MANISCHE EPISODEN
C2874871|T048||ICD10CM|MANIC EPISODE IN FULL REMISSION
C2874870|T048||ICD10CM|MANIC EPISODE IN PARTIAL REMISSION
C2874869|T048||ICD10CM|MANIC EPISODE, SEVERE WITH PSYCHOTIC SYMPTOMS
C2901789|T047|M86.069|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED TIBIA AND FIBULA|ACUTE HEMATOGENOUS OSTEOMYELITIS, UNSP TIBIA AND FIBULA
C2882342|T047|I63.111|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF RIGHT VERTEBRAL ARTERY|CEREBRAL INFARCTION DUE TO EMBOLISM OF R VERTEB ART
C2882343|T047|I63.112|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF LEFT VERTEBRAL ARTERY|CEREBRAL INFARCTION DUE TO EMBOLISM OF LEFT VERTEBRAL ARTERY
C4268477|T047|I63.113|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF BILATERAL VERTEBRAL ARTERIES|CEREBRAL INFARCTION DUE TO EMBOLISM OF BILATERAL VERTEB ART
C2901787|T047|M86.061|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, RIGHT TIBIA AND FIBULA|ACUTE HEMATOGENOUS OSTEOMYELITIS, RIGHT TIBIA AND FIBULA
C2859160|T037|S73.006A|ICD10CM|UNSPECIFIED DISLOCATION OF UNSPECIFIED HIP, INITIAL ENCOUNTER|UNSPECIFIED DISLOCATION OF UNSPECIFIED HIP, INIT ENCNTR
C2901788|T047|M86.062|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, LEFT TIBIA AND FIBULA|ACUTE HEMATOGENOUS OSTEOMYELITIS, LEFT TIBIA AND FIBULA
C2882344|T047|I63.119|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF UNSPECIFIED VERTEBRAL ARTERY|CEREBRAL INFARCTION DUE TO EMBOLISM OF UNSP VERTEBRAL ARTERY
C2833961|T037|S14.132D|ICD10CM|ANTERIOR CORD SYNDROME AT C2 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|ANTERIOR CORD SYNDROME AT C2, SUBS
C2833960|T037|S14.132A|ICD10CM|ANTERIOR CORD SYNDROME AT C2 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|ANTERIOR CORD SYNDROME AT C2, INIT
C2874259|T047|E72.09|ICD10CM|OTHER DISORDERS OF AMINO-ACID TRANSPORT|OTHER DISORDERS OF AMINO-ACID TRANSPORT
C2874803|T048|F19.180|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE ABUSE WITH PSYCHOACTIVE SUBSTANCE-INDUCED ANXIETY DISORDER|OTH PSYCHOACTIVE SUBSTANCE ABUSE W ANXIETY DISORDER
C0837058|T047|E13.00|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH HYPEROSMOLARITY WITHOUT NONKETOTIC HYPERGLYCEMIC-HYPEROSMOLAR COMA (NKHHC)|OTH DIAB W HYPROSM W/O NONKET HYPRGLY-HYPROS COMA (NKHHC)
C0837059|T047|E13.01|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH HYPEROSMOLARITY WITH COMA|OTH DIABETES MELLITUS WITH HYPEROSMOLARITY WITH COMA
C2833962|T037|S14.132S|ICD10CM|ANTERIOR CORD SYNDROME AT C2 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|ANTERIOR CORD SYNDROME AT C2, SEQUELA
C0340643|T046|I71.0|ICD10CM|DISSECTION OF UNSPECIFIED SITE OF AORTA|DISSECTION OF AORTA
C0340644|T047|I71.01|ICD10CM|DISSECTION OF THORACIC AORTA|DISSECTION OF THORACIC AORTA
C0837143|T047|I71.02|ICD10CM|DISSECTION OF ABDOMINAL AORTA|DISSECTION OF ABDOMINAL AORTA
C0837144|T047|I71.03|ICD10CM|DISSECTION OF THORACOABDOMINAL AORTA|DISSECTION OF THORACOABDOMINAL AORTA
C2905759|T037|X78.2XXD|ICD10CM|INTENTIONAL SELF-HARM BY SWORD OR DAGGER, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY SWORD OR DAGGER, SUBS ENCNTR
C0268548|T047|E72.21|ICD10CM|ARGININEMIA|ARGININEMIA
C0220994|T047|E72.20|ICD10CM|DISORDER OF UREA CYCLE METABOLISM, UNSPECIFIED|HYPERAMMONEMIA
C0175683|T047|E72.23|ICD10CM|CITRULLINEMIA|CITRULLINEMIA
C0596122|T046||ICD10CM|ARGINOSUCCINIC ACIDURIA
C2832064|T037|S06.302S|ICD10CM|UNSPECIFIED FOCAL TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|UNSP FOCAL TBI W LOSS OF CONSCIOUSNESS OF 31-59 MIN, SEQUELA
C2882388|T047|I63.429|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF UNSPECIFIED ANTERIOR CEREBRAL ARTERY|CEREBRAL INFRC DUE TO EMBOLISM OF UNSP ANT CEREBRAL ARTERY
C2874261|T047|E72.29|ICD10CM|OTHER DISORDERS OF UREA CYCLE METABOLISM|OTHER DISORDERS OF UREA CYCLE METABOLISM
C2890084|T037|T82.535A|ICD10CM|LEAKAGE OF UMBRELLA DEVICE, INITIAL ENCOUNTER|LEAKAGE OF UMBRELLA DEVICE, INITIAL ENCOUNTER
C2869759|T037|S98.012A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT FOOT AT ANKLE LEVEL, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMP OF LEFT FOOT AT ANKLE LEVEL, INIT
C2832590|T037|S06.820A|ICD10CM|INJURY OF LEFT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|INJURY OF L INT CAROTID, INTCR W/O LOC, INIT
C2833878|T037|S14.109A|ICD10CM|UNSPECIFIED INJURY AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY AT UNSP LEVEL OF CERVICAL SPINAL CORD, INIT
C0268641|T047|E72.00|ICD10CM|DISORDERS OF AMINO-ACID TRANSPORT, UNSPECIFIED|DISORDERS OF AMINO-ACID TRANSPORT, UNSPECIFIED
C2833879|T037|S14.109D|ICD10CM|UNSPECIFIED INJURY AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY AT UNSP LEVEL OF CERVICAL SPINAL CORD, SUBS
C4269263|T037|S02.111S|ICD10CM|TYPE II OCCIPITAL CONDYLE FRACTURE, UNSPECIFIED SIDE, SEQUELA|TYPE II OCCIPITAL CONDYLE FRACTURE, UNSP SIDE, SEQUELA
C2889228|T047|M05.379|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP ANK/FT
C2889226|T047|M05.371|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF RIGHT ANK/FT
C2889227|T047|M05.372|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF LEFT ANK/FT
C4269259|T037|S02.111B|ICD10CM|TYPE II OCCIPITAL CONDYLE FRACTURE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE II OCCIPITAL CONDYLE FRACTURE, UNSPECIFIED SIDE, 7THB
C4269258|T037|S02.111A|ICD10CM|TYPE II OCCIPITAL CONDYLE FRACTURE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE II OCCIPITAL CONDYLE FRACTURE, UNSPECIFIED SIDE, INIT
C2833168|T037|S12.030B|ICD10CM|DISPLACED POSTERIOR ARCH FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISPL POST ARCH FX FIRST CERVCAL VERTEBRA, INIT FOR OPN FX
C2874123|T047||ICD10CM|TYPE 2 DIABETES MELLITUS WITH HYPERGLYCEMIA
C2833167|T037|S12.030A|ICD10CM|DISPLACED POSTERIOR ARCH FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED POSTERIOR ARCH FX FIRST CERVCAL VERTEBRA, INIT
C0342262|T047|E11.69|ICD10AM|TYPE 2 DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATION|TYPE 2 DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATION
C2886161|T037|T65.822S|ICD10CM|TOXIC EFFECT OF HARMFUL ALGAE AND ALGAE TOXINS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFF OF HARMFUL ALGAE AND ALGAE TOXINS, SLF-HRM, SQLA
C2835398|T037|S22.069A|ICD10CM|UNSPECIFIED FRACTURE OF T7-T8 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF T7-T8 VERTEBRA, INIT FOR CLOS FX
C0432453|T047|Q95.3|DMDICD10|BALANCED SEX/AUTOSOMAL REARRANGEMENT IN ABNORMAL INDIVIDUAL|BALANCIERTES REARRANGEMENT ZWISCHEN GONOSOMEN UND AUTOSOMEN BEIM ABNORMEN INDIVIDUUM
C2856983|T037|S72.063B|ICD10CM|DISPLACED ARTICULAR FRACTURE OF HEAD OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL ARTIC FX HEAD OF UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2835399|T037|S22.069B|ICD10CM|UNSPECIFIED FRACTURE OF T7-T8 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF T7-T8 VERTEBRA, INIT FOR OPN FX
C2869838|T037|S98.212A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF TWO OR MORE LEFT LESSER TOES, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMP OF TWO OR MORE LEFT LESSER TOES, INIT
C2911407|T033|Z89.412|ICD10CM|ACQUIRED ABSENCE OF LEFT GREAT TOE|ACQUIRED ABSENCE OF LEFT GREAT TOE
C3264401|T047|J84.17|ICD10CM|OTHER INTERSTITIAL PULMONARY DISEASES WITH FIBROSIS IN DISEASES CLASSIFIED ELSEWHERE|OTH INTERSTIT PULMON DIS W FIBROSIS IN DIS CLASSD ELSWHR
C3264396|T047|J84.10|ICD10CM|PULMONARY FIBROSIS, UNSPECIFIED|PULMONARY FIBROSIS, UNSPECIFIED
C2890295|T037|T83.21XA|ICD10CM|BREAKDOWN (MECHANICAL) OF GRAFT OF URINARY ORGAN, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF GRAFT OF URINARY ORGAN, INIT
C2832598|T037|S06.822A|ICD10CM|INJURY OF LEFT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|INJURY OF L INT CAROTID, INTCR W LOC OF 31-59 MIN, INIT
C2901089|T046|M84.475A|ICD10CM|PATHOLOGICAL FRACTURE, LEFT FOOT, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, LEFT FOOT, INIT ENCNTR FOR FRACTURE
C2831616|T037|S02.92XB|ICD10CM|UNSPECIFIED FRACTURE OF FACIAL BONES, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF FACIAL BONES, INIT ENCNTR FOR OPEN FRACTURE
C2831615|T037|S02.92XA|ICD10CM|UNSPECIFIED FRACTURE OF FACIAL BONES, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF FACIAL BONES, INIT FOR CLOS FX
C2843329|T037|S48.919A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED SHOULDER AND UPPER ARM, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|COMPLETE TRAUM AMP OF UNSP SHLDR/UP ARM, LEVEL UNSP, INIT
C2833495|T037|S12.451B|ICD10CM|OTHER TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH TRAUM NONDISP SPONDYLOLYSIS OF 5TH CERVCAL VERT, 7THB
C2833494|T037|S12.451A|ICD10CM|OTHER TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH TRAUM NONDISP SPONDYLOLYSIS OF FIFTH CERVCAL VERT, INIT
C2831620|T037|S02.92XS|ICD10CM|UNSPECIFIED FRACTURE OF FACIAL BONES, SEQUELA|UNSPECIFIED FRACTURE OF FACIAL BONES, SEQUELA
C2843331|T037|S48.919S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED SHOULDER AND UPPER ARM, LEVEL UNSPECIFIED, SEQUELA|COMPLETE TRAUM AMP OF UNSP SHLDR/UP ARM, LEVEL UNSP, SEQUELA
C2865533|T037|S88.022A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT KNEE LEVEL, LEFT LOWER LEG, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION AT KNEE LEVEL, L LOW LEG, INIT
C2832391|T037|S06.381A|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF BRAINSTEM WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|CONTUS/LAC/HEM BRAINSTEM W LOC OF 30 MINUTES OR LESS, INIT
C2838680|T037|S34.124S|ICD10CM|INCOMPLETE LESION OF L4 LEVEL OF LUMBAR SPINAL CORD, SEQUELA|INCOMPLETE LESION OF L4 LEVEL OF LUMBAR SPINAL CORD, SEQUELA
C2874604|T048|F14.282|ICD10CM|COCAINE DEPENDENCE WITH COCAINE-INDUCED SLEEP DISORDER|COCAINE DEPENDENCE WITH COCAINE-INDUCED SLEEP DISORDER
C2874603|T048|F14.281|ICD10CM|COCAINE DEPENDENCE WITH COCAINE-INDUCED SEXUAL DYSFUNCTION|COCAINE DEPENDENCE WITH COCAINE-INDUCED SEXUAL DYSFUNCTION
C2900469|T047|A98.5|ICD10CM|HEMORRHAGIC FEVER WITH RENAL SYNDROME|SONGO FEVER
C2838679|T037|S34.124D|ICD10CM|INCOMPLETE LESION OF L4 LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|INCOMPLETE LESION OF L4 LEVEL OF LUMBAR SPINAL CORD, SUBS
C4268240|T048|F14.288|ICD10CM|COCAINE DEPENDENCE WITH OTHER COCAINE-INDUCED DISORDER|COCAINE USE DISORDER, SEVERE, WITH COCAINE-INDUCED OBSESSIVE COMPULSIVE OR RELATED DISORDER
C0155919|T047|J81.0|ICD10CM|ACUTE PULMONARY EDEMA|ACUTE PULMONARY EDEMA
C2832109|T037|S06.313S|ICD10CM|CONTUSION AND LACERATION OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, SEQUELA|CONTUS/LAC RIGHT CEREBRUM W LOC OF 1-5 HRS 59 MIN, SEQUELA
C2869773|T037|S98.022D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT FOOT AT ANKLE LEVEL, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMP OF LEFT FOOT AT ANKLE LEVEL, SUBS
C2977849|T037|S32.502B|ICD10CM|UNSPECIFIED FRACTURE OF LEFT PUBIS, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF LEFT PUBIS, INIT ENCNTR FOR OPEN FRACTURE
C0264694|T047|I25|DMDICD10|CHRONIC ISCHEMIC HEART DISEASE, UNSPECIFIED|CHRONISCHE ISCHAEMISCHE HERZKRANKHEIT
C0340291|T047|I25.6|DMDICD10|SILENT MYOCARDIAL ISCHEMIA|STUMME MYOKARDISCHAEMIE
C2837713|T037|S32.122A|ICD10CM|SEVERELY DISPLACED ZONE II FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SEVERELY DISPLACED ZONE II FRACTURE OF SACRUM, INIT
C2832107|T037|S06.313A|ICD10CM|CONTUSION AND LACERATION OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|CONTUS/LAC RIGHT CEREBRUM W LOC OF 1-5 HRS 59 MIN, INIT
C0349782|T047|I25.5|DMDICD10|ISCHEMIC CARDIOMYOPATHY|ISCHAEMISCHE KARDIOMYOPATHIE
C2882169|T046|I25.2|ICD10CM|OLD MYOCARDIAL INFARCTION|PAST MYOCARDIAL INFARCTION DIAGNOSED BY ECG OR OTHER INVESTIGATION, BUT CURRENTLY PRESENTING NO SYMPTOMS
C1541919|T047||ICD10CM|ANEURYSM OF HEART
C2845943|T191|C74.10|ICD10CM|MALIGNANT NEOPLASM OF MEDULLA OF UNSPECIFIED ADRENAL GLAND|MALIGNANT NEOPLASM OF MEDULLA OF UNSPECIFIED ADRENAL GLAND
C2845944|T191|C74.11|ICD10CM|MALIGNANT NEOPLASM OF MEDULLA OF RIGHT ADRENAL GLAND|MALIGNANT NEOPLASM OF MEDULLA OF RIGHT ADRENAL GLAND
C2845945|T191|C74.12|ICD10CM|MALIGNANT NEOPLASM OF MEDULLA OF LEFT ADRENAL GLAND|MALIGNANT NEOPLASM OF MEDULLA OF LEFT ADRENAL GLAND
C2878845|T037|T44.4X2S|ICD10CM|POISONING BY PREDOMINANTLY ALPHA-ADRENORECEPTOR AGONISTS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY PREDOM ALPHA-ADRENOCPT AGONISTS, SELF-HARM, SEQUELA
C2876166|T037|T31.83|ICD10CM|BURNS INVOLVING 80-89% OF BODY SURFACE WITH 30-39% THIRD DEGREE BURNS|BURNS OF 80-89% OF BODY SURFACE W 30-39% THIRD DEGREE BURNS
C2876165|T037|T31.82|ICD10CM|BURNS INVOLVING 80-89% OF BODY SURFACE WITH 20-29% THIRD DEGREE BURNS|BURNS OF 80-89% OF BODY SURFACE W 20-29% THIRD DEGREE BURNS
C2878843|T037|T44.4X2A|ICD10CM|POISONING BY PREDOMINANTLY ALPHA-ADRENORECEPTOR AGONISTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY PREDOM ALPHA-ADRENOCPT AGONISTS, SELF-HARM, INIT
C1264197|T191|C09.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF TONSIL|BOESARTIGE NEUBILDUNG: TONSILLE, MEHRERE TEILBEREICHE UEBERLAPPEND
C1719638|T046||ICD10CM|UNSPECIFIED CONVULSIONS
C2845929|T191|C72.20|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED OLFACTORY NERVE|MALIGNANT NEOPLASM OF UNSPECIFIED OLFACTORY NERVE
C4267950|T047|E08.37X1|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, RIGHT EYE|DIAB WITH DIABETIC MACULAR EDEMA, RESOLVED FOL TRTMT, R EYE
C4267951|T047|E08.37X2|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, LEFT EYE|DIAB WITH DIAB MACULAR EDEMA, RESOLVED FOL TRTMT, LEFT EYE
C4267952|T047|E08.37X3|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, BILATERAL|DIABETES WITH DIABETIC MACULAR EDEMA, RESOLVED FOL TRTMT, BI
C2921125|T047|R56.1|ICD10CM|POST TRAUMATIC SEIZURES|POST TRAUMATIC SEIZURES
C2865535|T037|S88.022S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT KNEE LEVEL, LEFT LOWER LEG, SEQUELA|PARTIAL TRAUMATIC AMP AT KNEE LEVEL, L LOW LEG, SEQUELA
C4267953|T047|E08.37X9|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, UNSPECIFIED EYE|DIAB WITH DIABETIC MACULAR EDEMA, RESOLVED FOL TRTMT, UNSP
C2853992|T191|C84.91|ICD10CM|MATURE T/NK-CELL LYMPHOMAS, UNSPECIFIED, LYMPH NODES OF HEAD, FACE, AND NECK|MATURE T/NK-CELL LYMPH, UNSP, NODES OF HEAD, FACE, AND NECK
C2853991|T191|C84.90|ICD10CM|MATURE T/NK-CELL LYMPHOMAS, UNSPECIFIED, UNSPECIFIED SITE|MATURE T/NK-CELL LYMPHOMAS, UNSPECIFIED, UNSPECIFIED SITE
C2853994|T191|C84.93|ICD10CM|MATURE T/NK-CELL LYMPHOMAS, UNSPECIFIED, INTRA-ABDOMINAL LYMPH NODES|MATURE T/NK-CELL LYMPHOMAS, UNSP, INTRA-ABD LYMPH NODES
C2853993|T191|C84.92|ICD10CM|MATURE T/NK-CELL LYMPHOMAS, UNSPECIFIED, INTRATHORACIC LYMPH NODES|MATURE T/NK-CELL LYMPHOMAS, UNSP, INTRATHORACIC LYMPH NODES
C2853996|T191|C84.95|ICD10CM|MATURE T/NK-CELL LYMPHOMAS, UNSPECIFIED, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|MATURE T/NK-CELL LYMPH, UNSP, NODES OF ING RGN AND LOW LIMB
C2889404|T047|M06.059|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, UNSPECIFIED HIP|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, UNSP HIP
C2853998|T191|C84.97|ICD10CM|MATURE T/NK-CELL LYMPHOMAS, UNSPECIFIED, SPLEEN|MATURE T/NK-CELL LYMPHOMAS, UNSPECIFIED, SPLEEN
C2853997|T191|C84.96|ICD10CM|MATURE T/NK-CELL LYMPHOMAS, UNSPECIFIED, INTRAPELVIC LYMPH NODES|MATURE T/NK-CELL LYMPHOMAS, UNSP, INTRAPELVIC LYMPH NODES
C2854000|T191|C84.99|ICD10CM|MATURE T/NK-CELL LYMPHOMAS, UNSPECIFIED, EXTRANODAL AND SOLID ORGAN SITES|MATURE T/NK-CELL LYMPH, UNSP, EXTRNOD AND SOLID ORGAN SITES
C2853999|T191|C84.98|ICD10CM|MATURE T/NK-CELL LYMPHOMAS, UNSPECIFIED, LYMPH NODES OF MULTIPLE SITES|MATURE T/NK-CELL LYMPHOMAS, UNSP, LYMPH NODES MULT SITE
C4267947|T047|E08.3593|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|DIAB WITH PROLIF DIABETIC RTNOP WITHOUT MACULAR EDEMA, BI
C4267946|T047|E08.3592|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|DIAB WITH PROLIF DIAB RTNOP WITHOUT MACULAR EDEMA, LEFT EYE
C2902379|T047|M89.671|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, RIGHT ANKLE AND FOOT|OSTEOPATHY AFTER POLIOMYELITIS, RIGHT ANKLE AND FOOT
C2889402|T047|M06.051|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, RIGHT HIP|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, RIGHT HIP
C2889403|T047|M06.052|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, LEFT HIP|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, LEFT HIP
C2902380|T047|M89.672|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, LEFT ANKLE AND FOOT|OSTEOPATHY AFTER POLIOMYELITIS, LEFT ANKLE AND FOOT
C2835168|T037|S22.002A|ICD10CM|UNSTABLE BURST FRACTURE OF UNSPECIFIED THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSTABLE BURST FRACTURE OF UNSP THORACIC VERTEBRA, INIT
C2869863|T037|S98.311S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT MIDFOOT, SEQUELA|COMPLETE TRAUMATIC AMPUTATION OF RIGHT MIDFOOT, SEQUELA
C2869862|T037|S98.311D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT MIDFOOT, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF RIGHT MIDFOOT, SUBS ENCNTR
C0864957|T191|C51.9|ICD10CM|MALIGNANT NEOPLASM OF VULVA, UNSPECIFIED|MALIGNANT NEOPLASM OF PUDENDUM
C1263790|T191|C51.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF VULVA|BOESARTIGE NEUBILDUNG: VULVA, MEHRERE TEILBEREICHE UEBERLAPPEND
C2869861|T037|S98.311A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT MIDFOOT, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF RIGHT MIDFOOT, INIT ENCNTR
C0153589|T191|C51.2|DMDICD10|MALIGNANT NEOPLASM OF CLITORIS|BOESARTIGE NEUBILDUNG DER VULVA: KLITORIS
C0496815|T191|C51.1|DMDICD10|MALIGNANT NEOPLASM OF LABIUM MINUS|BOESARTIGE NEUBILDUNG DER VULVA: LABIUM MINUS
C2842144|T191|C51.0|ICD10CM|MALIGNANT NEOPLASM OF LABIUM MAJUS|MALIGNANT NEOPLASM OF BARTHOLIN'S [GREATER VESTIBULAR] GLAND
C2869853|T037|S98.222S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF TWO OR MORE LEFT LESSER TOES, SEQUELA|PARTIAL TRAUM AMP OF TWO OR MORE LEFT LESSER TOES, SEQUELA
C3161074|T046|D61.811|ICD10CM|OTHER DRUG-INDUCED PANCYTOPENIA|OTHER DRUG-INDUCED PANCYTOPENIA
C2869852|T037|S98.222D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF TWO OR MORE LEFT LESSER TOES, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMP OF TWO OR MORE LEFT LESSER TOES, SUBS
C2869851|T037|S98.222A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF TWO OR MORE LEFT LESSER TOES, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP OF TWO OR MORE LEFT LESSER TOES, INIT
C0694477|T047|G63|DMDICD10|POLYNEUROPATHY IN DISEASES CLASSIFIED ELSEWHERE|POLYNEUROPATHIE BEI ANDERENORTS KLASSIFIZIERTEN KRANKHEITEN
C0477401|T047|G64|DMDICD10|OTHER DISORDERS OF PERIPHERAL NERVOUS SYSTEM|SONSTIGE KRANKHEITEN DES PERIPHEREN NERVENSYSTEMS
C2895184|T047|M33.11|ICD10CM|OTHER DERMATOMYOSITIS WITH RESPIRATORY INVOLVEMENT|OTHER DERMATOMYOSITIS WITH RESPIRATORY INVOLVEMENT
C4509351|T047|M33.10|ICD10CM|OTHER DERMATOMYOSITIS, ORGAN INVOLVEMENT UNSPECIFIED|OTHER DERMATOMYOSITIS, ORGAN INVOLVEMENT UNSPECIFIED
C4509352|T047|M33.13|ICD10CM|OTHER DERMATOMYOSITIS WITHOUT MYOPATHY|OTHER DERMATOMYOSITIS WITHOUT MYOPATHY
C2895185|T047|M33.12|ICD10CM|OTHER DERMATOMYOSITIS WITH MYOPATHY|OTHER DERMATOMYOSITIS WITH MYOPATHY
C4270359|T046|T83.62XA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO IMPLANTED TESTICULAR PROSTHESIS, INITIAL ENCOUNTER|I/I REACT D/T IMPLANTED TESTICULAR PROSTHESIS, INIT
C4509353|T047|M33.19|ICD10CM|OTHER DERMATOMYOSITIS WITH OTHER ORGAN INVOLVEMENT|OTHER DERMATOMYOSITIS WITH OTHER ORGAN INVOLVEMENT
C2832278|T037|S06.354A|ICD10CM|TRAUMATIC HEMORRHAGE OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|TRAUM HEMOR LEFT CEREBRUM W LOC OF 6 HOURS TO 24 HOURS, INIT
C2858921|T037|S72.465C|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP SUPRCNDL FX W INTRCNDL EXTN LOW END L FEMR, 7THC
C2857344|T037|S72.126C|ICD10CM|NONDISPLACED FRACTURE OF LESSER TROCHANTER OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF LESS TROCHANTER OF UNSP FEMR, 7THC
C2882206|T047|I25.798|ICD10CM|ATHEROSCLEROSIS OF OTHER CORONARY ARTERY BYPASS GRAFT(S) WITH OTHER FORMS OF ANGINA PECTORIS|ATHEROSCLEROSIS OF CABG W OTH ANGINA PECTORIS
C2882207|T047|I25.799|ICD10CM|ATHEROSCLEROSIS OF OTHER CORONARY ARTERY BYPASS GRAFT(S) WITH UNSPECIFIED ANGINA PECTORIS|ATHEROSCLEROSIS OF CABG W UNSP ANGINA PECTORIS
C2832280|T037|S06.354S|ICD10CM|TRAUMATIC HEMORRHAGE OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|TRAUM HEMOR LEFT CEREBRUM W LOC OF 6-24 HRS, SEQUELA
C2882204|T047|I25.790|ICD10CM|ATHEROSCLEROSIS OF OTHER CORONARY ARTERY BYPASS GRAFT(S) WITH UNSTABLE ANGINA PECTORIS|ATHEROSCLEROSIS OF CABG W UNSTABLE ANGINA PECTORIS
C2882205|T047|I25.791|ICD10CM|ATHEROSCLEROSIS OF OTHER CORONARY ARTERY BYPASS GRAFT(S) WITH ANGINA PECTORIS WITH DOCUMENTED SPASM|ATHEROSCLEROSIS OF CABG W ANGINA PECTORIS W DOCUMENTED SPASM
C2853822|T191|C82.35|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|FOLICLAR LYMPH GRADE IIIA, NODES OF ING RGN AND LOWER LIMB
C2853821|T191|C82.34|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIA, LYMPH NODES OF AXILLA AND UPPER LIMB|FOLICLAR LYMPHOMA GRADE IIIA, NODES OF AXILLA AND UPPER LIMB
C2853824|T191|C82.37|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIA, SPLEEN|FOLLICULAR LYMPHOMA GRADE IIIA, SPLEEN
C2853823|T191|C82.36|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIA, INTRAPELVIC LYMPH NODES|FOLLICULAR LYMPHOMA GRADE IIIA, INTRAPELVIC LYMPH NODES
C2853818|T191|C82.31|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIA, LYMPH NODES OF HEAD, FACE, AND NECK|FOLICLAR LYMPHOMA GRADE IIIA, NODES OF HEAD, FACE, AND NECK
C2853817|T191|C82.30|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIA, UNSPECIFIED SITE|FOLLICULAR LYMPHOMA GRADE IIIA, UNSPECIFIED SITE
C2853820|T191|C82.33|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIA, INTRA-ABDOMINAL LYMPH NODES|FOLLICULAR LYMPHOMA GRADE IIIA, INTRA-ABDOMINAL LYMPH NODES
C2853819|T191|C82.32|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIA, INTRATHORACIC LYMPH NODES|FOLLICULAR LYMPHOMA GRADE IIIA, INTRATHORACIC LYMPH NODES
C2882678|T046|I69.963|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING RIGHT NON-DOMINANT SIDE|OTH PARLYT SYND FOL UNSP CEREBVASC DIS AFF RIGHT NONDOM SIDE
C2882369|T047|I63.322|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF LEFT ANTERIOR CEREBRAL ARTERY|CEREBRAL INFRC DUE TO THOMBOS OF LEFT ANT CEREBRAL ARTERY
C2882676|T046|I69.961|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING RIGHT DOMINANT SIDE|OTH PARLYT SYND FOL UNSP CEREBVASC DIS AFF RIGHT DOM SIDE
C2873894|T047|E08.29|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH OTHER DIABETIC KIDNEY COMPLICATION|DIABETES DUE TO UNDRL CONDITION W OTH DIABETIC KIDNEY COMP
C2853826|T191|C82.39|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIA, EXTRANODAL AND SOLID ORGAN SITES|FOLICLAR LYMPHOMA GRADE IIIA, EXTRNOD AND SOLID ORGAN SITES
C2853825|T191|C82.38|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIA, LYMPH NODES OF MULTIPLE SITES|FOLLICULAR LYMPHOMA GRADE IIIA, LYMPH NODES MULT SITE
C2882680|T046|I69.965|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE, BILATERAL|OTH PARALYTIC SYNDROME FOLLOWING UNSP CEREBVASC DISEASE, BI
C2882679|T046|I69.964|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING LEFT NON-DOMINANT SIDE|OTH PARLYT SYND FOL UNSP CEREBVASC DIS AFF LEFT NONDOM SIDE
C0030807|T047|L10|DMDICD10|PEMPHIGUS, UNSPECIFIED|PEMPHIGUSKRANKHEITEN
C2835313|T037|S22.042B|ICD10CM|UNSTABLE BURST FRACTURE OF FOURTH THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSTABLE BURST FX FOURTH THOR VERTEBRA, INIT FOR OPN FX
C2878635|T037|T43.632A|ICD10CM|POISONING BY METHYLPHENIDATE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY METHYLPHENIDATE, INTENTIONAL SELF-HARM, INIT
C0263316|T047|L10.1|DMDICD10|PEMPHIGUS VEGETANS|PEMPHIGUS VEGETANS
C0030809|T047|L10.0|DMDICD10|PEMPHIGUS VULGARIS|PEMPHIGUS VULGARIS
C0263314|T047|L10.3|DMDICD10|BRAZILIAN PEMPHIGUS [FOGO SELVAGEM]|BRASILIANISCHER PEMPHIGUS [FOGO SELVAGEM]
C0263313|T047|L10.2|DMDICD10|PEMPHIGUS FOLIACEOUS|PEMPHIGUS FOLIACEUS
C0451938|T046|L10.5|DMDICD10|DRUG-INDUCED PEMPHIGUS|ARZNEIMITTELINDUZIERTER PEMPHIGUS
C0263312|T047|L10.4|DMDICD10|PEMPHIGUS ERYTHEMATOSUS|PEMPHIGUS ERYTHEMATOSUS
C2887226|T047|I83.224|ICD10CM|VARICOSE VEINS OF LEFT LOWER EXTREMITY WITH BOTH ULCER OF HEEL AND MIDFOOT AND INFLAMMATION|VARICOS VN OF L LOW EXTREM W ULC OF HEEL & MIDFT AND INFLAM
C2887228|T047|I83.225|ICD10CM|VARICOSE VEINS OF LEFT LOWER EXTREMITY WITH BOTH ULCER OTHER PART OF FOOT AND INFLAMMATION|VARICOS VN OF L LOW EXTREM W ULC OTH PART OF FOOT AND INFLAM
C4269476|T037|S02.622B|ICD10CM|FRACTURE OF SUBCONDYLAR PROCESS OF LEFT MANDIBLE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF SUBCONDYLAR PROCESS OF LEFT MANDIBLE, 7THB
C2887222|T047|I83.221|ICD10CM|VARICOSE VEINS OF LEFT LOWER EXTREMITY WITH BOTH ULCER OF THIGH AND INFLAMMATION|VARICOS VN OF L LOW EXTREM W ULC OF THIGH AND INFLAMMATION
C2887223|T047|I83.222|ICD10CM|VARICOSE VEINS OF LEFT LOWER EXTREMITY WITH BOTH ULCER OF CALF AND INFLAMMATION|VARICOS VN OF L LOW EXTREM W ULC OF CALF AND INFLAMMATION
C2887224|T047|I83.223|ICD10CM|VARICOSE VEINS OF LEFT LOWER EXTREMITY WITH BOTH ULCER OF ANKLE AND INFLAMMATION|VARICOS VN OF L LOW EXTREM W ULC OF ANKLE AND INFLAMMATION
C2887229|T047|I83.228|ICD10CM|VARICOSE VEINS OF LEFT LOWER EXTREMITY WITH BOTH ULCER OF OTHER PART OF LOWER EXTREMITY AND INFLAMMATION|VARICOS VN OF L LOW EXTREM W ULC OTH PRT LOW EXTRM & INFLAM
C2887230|T047|I83.229|ICD10CM|VARICOSE VEINS OF LEFT LOWER EXTREMITY WITH BOTH ULCER OF UNSPECIFIED SITE AND INFLAMMATION|VARICOS VN OF L LOW EXTREM W ULC OF UNSP SITE AND INFLAM
C4269480|T037|S02.622S|ICD10CM|FRACTURE OF SUBCONDYLAR PROCESS OF LEFT MANDIBLE, SEQUELA|FRACTURE OF SUBCONDYLAR PROCESS OF LEFT MANDIBLE, SEQUELA
C2890750|T037|T84.318A|ICD10CM|BREAKDOWN (MECHANICAL) OF OTHER BONE DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|BREAKDOWN OF BONE DEVICES, IMPLANTS AND GRAFTS, INIT
C2885509|T037|T63.2X2S|ICD10CM|TOXIC EFFECT OF VENOM OF SCORPION, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF SCORPION, SELF-HARM, SEQUELA
C2837626|T037|S32.050B|ICD10CM|WEDGE COMPRESSION FRACTURE OF FIFTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|WEDGE COMPRSN FX FIFTH LUM VERTEBRA, INIT FOR OPN FX
C2837625|T037|S32.050A|ICD10CM|WEDGE COMPRESSION FRACTURE OF FIFTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|WEDGE COMPRESSION FRACTURE OF FIFTH LUMBAR VERTEBRA, INIT
C2885237|T037|T62.1X2A|ICD10CM|TOXIC EFFECT OF INGESTED BERRIES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF INGESTED BERRIES, SELF-HARM, INIT
C2901839|T047|M86.279|ICD10CM|SUBACUTE OSTEOMYELITIS, UNSPECIFIED ANKLE AND FOOT|SUBACUTE OSTEOMYELITIS, UNSPECIFIED ANKLE AND FOOT
C2901837|T047|M86.271|ICD10CM|SUBACUTE OSTEOMYELITIS, RIGHT ANKLE AND FOOT|SUBACUTE OSTEOMYELITIS, RIGHT ANKLE AND FOOT
C2901838|T047|M86.272|ICD10CM|SUBACUTE OSTEOMYELITIS, LEFT ANKLE AND FOOT|SUBACUTE OSTEOMYELITIS, LEFT ANKLE AND FOOT
C2831935|T037|S06.0X0S|ICD10CM|CONCUSSION WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|CONCUSSION WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA
C2890770|T037|T84.398A|ICD10CM|OTHER MECHANICAL COMPLICATION OF OTHER BONE DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|MECH COMPL OF OTH BONE DEVICES, IMPLANTS AND GRAFTS, INIT
C2875180|T047|G43.809|ICD10CM|OTHER MIGRAINE, NOT INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|OTHER MIGRAINE, NOT INTRACTABLE, WITHOUT STATUS MIGRAINOSUS
C2831974|T037|S06.1X0S|ICD10CM|TRAUMATIC CEREBRAL EDEMA WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|TRAUMATIC CEREBRAL EDEMA W/O LOSS OF CONSCIOUSNESS, SEQUELA
C2875179|T047|G43.801|ICD10CM|OTHER MIGRAINE, NOT INTRACTABLE, WITH STATUS MIGRAINOSUS|OTHER MIGRAINE, NOT INTRACTABLE, WITH STATUS MIGRAINOSUS
C2831972|T037|S06.1X0A|ICD10CM|TRAUMATIC CEREBRAL EDEMA WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|TRAUMATIC CEREBRAL EDEMA W/O LOSS OF CONSCIOUSNESS, INIT
C2842034|T191|C47.22|ICD10CM|MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF LEFT LOWER LIMB, INCLUDING HIP|MALIG NEOPLASM OF PRPH NERVES OF LEFT LOWER LIMB, INC HIP
C2842033|T191|C47.21|ICD10CM|MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF RIGHT LOWER LIMB, INCLUDING HIP|MALIG NEOPLASM OF PRPH NERVES OF RIGHT LOWER LIMB, INC HIP
C2842032|T191|C47.20|ICD10CM|MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF UNSPECIFIED LOWER LIMB, INCLUDING HIP|MALIG NEOPLASM OF PRPH NERVES OF UNSP LOWER LIMB, INC HIP
C2833900|T037|S14.115S|ICD10CM|COMPLETE LESION AT C5 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|COMPLETE LESION AT C5 LEVEL OF CERVICAL SPINAL CORD, SEQUELA
C4509214|T047|I27.24|ICD10CM|CHRONIC THROMBOEMBOLIC PULMONARY HYPERTENSION|GROUP 4 PULMONARY HYPERTENSION
C4509213|T047|I27.23|ICD10CM|PULMONARY HYPERTENSION DUE TO LUNG DISEASES AND HYPOXIA|GROUP 3 PULMONARY HYPERTENSION
C4509211|T047|I27.22|ICD10CM|PULMONARY HYPERTENSION DUE TO LEFT HEART DISEASE|GROUP 2 PULMONARY HYPERTENSION
C4509210|T047|I27.21|ICD10CM|SECONDARY PULMONARY ARTERIAL HYPERTENSION|(ASSOCIATED) (DRUG-INDUCED) (TOXIN-INDUCED) (SECONDARY) GROUP 1 PULMONARY HYPERTENSION
C4509208|T047|I27.20|ICD10CM|PULMONARY HYPERTENSION, UNSPECIFIED|PULMONARY HYPERTENSION, UNSPECIFIED
C2833898|T037|S14.115A|ICD10CM|COMPLETE LESION AT C5 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION AT C5 LEVEL OF CERVICAL SPINAL CORD, INIT
C4509219|T047|I27.29|ICD10CM|OTHER SECONDARY PULMONARY HYPERTENSION|PULMONARY HYPERTENSION DUE TO OTHER SYSTEMIC DISORDERS
C2889589|T047|M08.452|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, LEFT HIP|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, LEFT HIP
C2885255|T037|T62.2X2S|ICD10CM|TOXIC EFFECT OF OTHER INGESTED (PARTS OF) PLANT(S), INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF INGEST (PARTS OF) PLANT(S), SLF-HRM, SEQUELA
C2889588|T047|M08.451|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, RIGHT HIP|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, RIGHT HIP
C2895343|T037|M48.58XA|ICD10CM|COLLAPSED VERTEBRA, NOT ELSEWHERE CLASSIFIED, SACRAL AND SACROCOCCYGEAL REGION, INITIAL ENCOUNTER FOR FRACTURE|COLLAPSED VERTEBRA, NEC, SACR/SACROCYGL REGION, INIT
C2861669|T191|D03.21|ICD10CM|MELANOMA IN SITU OF RIGHT EAR AND EXTERNAL AURICULAR CANAL|MELANOMA IN SITU OF RIGHT EAR AND EXTERNAL AURICULAR CANAL
C2889590|T047|M08.45|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED HIP|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, HIP
C2349872|T033|Z91.15|ICD10CM|PATIENT'S NONCOMPLIANCE WITH RENAL DIALYSIS|PATIENT'S NONCOMPLIANCE WITH RENAL DIALYSIS
C2856878|T037|S72.046A|ICD10CM|NONDISPLACED FRACTURE OF BASE OF NECK OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF BASE OF NECK OF UNSP FEMUR, INIT FOR CLOS FX
C2857223|T037|S72.115B|ICD10CM|NONDISPLACED FRACTURE OF GREATER TROCHANTER OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF GREATER TROCHANTER OF L FEMR, 7THB
C2856880|T037|S72.046C|ICD10CM|NONDISPLACED FRACTURE OF BASE OF NECK OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF BASE OF NK OF UNSP FEMR, 7THC
C2856879|T037|S72.046B|ICD10CM|NONDISPLACED FRACTURE OF BASE OF NECK OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF BASE OF NK OF UNSP FEMR, 7THB
C2835794|T037|S24.119S|ICD10CM|COMPLETE LESION AT UNSPECIFIED LEVEL OF THORACIC SPINAL CORD, SEQUELA|COMPLETE LESION AT UNSP LEVEL OF THOR SPINAL CORD, SEQUELA
C0268124|T047|D81.3|DMDICD10|ADENOSINE DEAMINASE [ADA] DEFICIENCY|ADENOSINDESAMINASE[ADA]-MANGEL
C0451694|T047|D81.2|DMDICD10|SEVERE COMBINED IMMUNODEFICIENCY [SCID] WITH LOW OR NORMAL B-CELL NUMBERS|SCHWERER KOMBINIERTER IMMUNDEFEKT [SCID] MIT NIEDRIGER ODER NORMALER B-ZELLEN-ZAHL
C0451693|T047|D81.1|DMDICD10|SEVERE COMBINED IMMUNODEFICIENCY [SCID] WITH LOW T- AND B-CELL NUMBERS|SCHWERER KOMBINIERTER IMMUNDEFEKT [SCID] MIT NIEDRIGER T- UND B-ZELLEN-ZAHL
C2531305|T061|D810|ICD10PCS|SEVERE COMBINED IMMUNODEFICIENCY [SCID] WITH RETICULAR DYSGENESIS|RADIATION THERAPY @ EYE @ BRACHYTHERAPY @ EYE
C0451696|T047|D81.7|DMDICD10|MAJOR HISTOCOMPATIBILITY COMPLEX CLASS II DEFICIENCY|HAUPTHISTOKOMPATIBILITAETS-KOMPLEX-KLASSE-II-DEFEKT [MHC-KLASSE-II-DEFEKT]
C0451695|T047|D81.6|DMDICD10|MAJOR HISTOCOMPATIBILITY COMPLEX CLASS I DEFICIENCY|HAUPTHISTOKOMPATIBILITAETS-KOMPLEX-KLASSE-I-DEFEKT [MHC-KLASSE-I-DEFEKT]
C0268125|T047|D81.5|DMDICD10|PURINE NUCLEOSIDE PHOSPHORYLASE [PNP] DEFICIENCY|PURINNUKLEOSID-PHOSPHORYLASE[PNP]-MANGEL
C0152094|T047|D81.4|DMDICD10|NEZELOF'S SYNDROME|NEZELOF-SYNDROM
C2873846|T047|D81.9|ICD10CM|COMBINED IMMUNODEFICIENCY, UNSPECIFIED|SEVERE COMBINED IMMUNODEFICIENCY DISORDER [SCID] NOS
C2835793|T037|S24.119D|ICD10CM|COMPLETE LESION AT UNSPECIFIED LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION AT UNSP LEVEL OF THORACIC SPINAL CORD, SUBS
C2857925|T037|S72.341A|ICD10CM|DISPLACED SPIRAL FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED SPIRAL FRACTURE OF SHAFT OF RIGHT FEMUR, INIT
C2835792|T037|S24.119A|ICD10CM|COMPLETE LESION AT UNSPECIFIED LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION AT UNSP LEVEL OF THORACIC SPINAL CORD, INIT
C2857926|T037|S72.341B|ICD10CM|DISPLACED SPIRAL FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL SPIRAL FX SHAFT OF R FEMUR, INIT FOR OPN FX TYPE I/2
C2884052|T037|T51.8X2A|ICD10CM|TOXIC EFFECT OF OTHER ALCOHOLS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF OTH ALCOHOLS, INTENTIONAL SELF-HARM, INIT
C2876818|T037|T37.1X2A|ICD10CM|POISONING BY ANTIMYCOBACTERIAL DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ANTIMYCOBACTERIAL DRUGS, SELF-HARM, INIT
C4268634|T047|K55.062|ICD10CM|DIFFUSE ACUTE INFARCTION OF INTESTINE, PART UNSPECIFIED|DIFFUSE ACUTE INFARCTION OF INTESTINE, PART UNSPECIFIED
C4268633|T047|K55.061|ICD10CM|FOCAL (SEGMENTAL) ACUTE INFARCTION OF INTESTINE, PART UNSPECIFIED|FOCAL ACUTE INFARCTION OF INTESTINE, PART UNSPECIFIED
C2896544|T046|M80.039A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, UNSPECIFIED FOREARM, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, UNSP FOREARM, INIT
C4268635|T047|K55.069|ICD10CM|ACUTE INFARCTION OF INTESTINE, PART AND EXTENT UNSPECIFIED|ACUTE INFARCTION OF INTESTINE, PART AND EXTENT UNSPECIFIED
C2890703|T037|T84.216A|ICD10CM|BREAKDOWN (MECHANICAL) OF INTERNAL FIXATION DEVICE OF VERTEBRAE, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF INT FIX OF VERTEBRAE, INIT
C2873816|T047|D72.0|ICD10CM|GENETIC ANOMALIES OF LEUKOCYTES|PELGER-HUËT (GRANULATION) (GRANULOCYTE) ANOMALY
C4267973|T047|E09.3419|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|DRUG/CHEM DIAB WITH SEVERE NONP RTNOP WITH MCLR EDEMA, UNSP
C2833973|T037|S14.135D|ICD10CM|ANTERIOR CORD SYNDROME AT C5 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|ANTERIOR CORD SYNDROME AT C5, SUBS
C4267970|T047|E09.3411|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|DRUG/CHEM DIAB WITH SEVERE NONP RTNOP WITH MCLR EDEMA, R EYE
C4267972|T047|E09.3413|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|DRUG/CHEM DIAB WITH SEVERE NONP RTNOP WITH MACULAR EDEMA, BI
C4267971|T047|E09.3412|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|DRUG/CHEM DIAB WITH SEVERE NONP RTNOP WITH MCLR EDEMA, L EYE
C2838632|T037|S34.105A|ICD10CM|UNSPECIFIED INJURY TO L5 LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY TO L5 LEVEL OF LUMBAR SPINAL CORD, INIT ENCNTR
C2860018|T037|S78.129A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN UNSPECIFIED HIP AND KNEE, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP AT LEVEL BETW UNSP HIP AND KNEE, INIT
C2838633|T037|S34.105D|ICD10CM|UNSPECIFIED INJURY TO L5 LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY TO L5 LEVEL OF LUMBAR SPINAL CORD, SUBS ENCNTR
C2860019|T037|S78.129D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN UNSPECIFIED HIP AND KNEE, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMP AT LEVEL BETW UNSP HIP AND KNEE, SUBS
C2887861|T047|K56.2|ICD10CM|VOLVULUS|TWIST OF COLON OR INTESTINE
C0156156|T047|K56.3|DMDICD10|GALLSTONE ILEUS|GALLENSTEINILEUS
C0267474|T047|K56.0|ICD10CM|PARALYTIC ILEUS|PARALYSIS OF COLON
C2887858|T046|K56.1|ICD10CM|INTUSSUSCEPTION|INTUSSUSCEPTION OR INVAGINATION OF RECTUM
C0348744|T047|K56.7|DMDICD10|ILEUS, UNSPECIFIED|ILEUS, NICHT NAEHER BEZEICHNET
C4509255|T047|K56.5|ICD10CM|INTESTINAL ADHESIONS [BANDS] WITH OBSTRUCTION (POSTPROCEDURAL) (POSTINFECTION)|PERITONEAL ADHESIONS [BANDS] WITH INTESTINAL OBSTRUCTION (POSTINFECTION)
C2860020|T037|S78.129S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN UNSPECIFIED HIP AND KNEE, SEQUELA|PARTIAL TRAUM AMP AT LEVEL BETW UNSP HIP AND KNEE, SEQUELA
C2889150|T047|M05.142|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT HAND|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT HAND
C2889149|T047|M05.141|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT HAND|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889306|T047|M05.631|ICD10CM|RHEUMATOID ARTHRITIS OF RIGHT WRIST WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF R WRIST W INVOLV OF ORGANS AND SYSTEMS
C2889307|T047|M05.632|ICD10CM|RHEUMATOID ARTHRITIS OF LEFT WRIST WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF L WRIST W INVOLV OF ORGANS AND SYSTEMS
C2889151|T047|M05.149|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP HAND
C2889308|T047|M05.639|ICD10CM|RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF UNSP WRIST W INVOLV OF ORGANS AND SYSTEMS
C2842058|T191|C4A.30|ICD10CM|MERKEL CELL CARCINOMA OF UNSPECIFIED PART OF FACE|MERKEL CELL CARCINOMA OF UNSPECIFIED PART OF FACE
C2842059|T191|C4A.31|ICD10CM|MERKEL CELL CARCINOMA OF NOSE|MERKEL CELL CARCINOMA OF NOSE
C2842060|T191|C4A.39|ICD10CM|MERKEL CELL CARCINOMA OF OTHER PARTS OF FACE|MERKEL CELL CARCINOMA OF OTHER PARTS OF FACE
C0018197|T191|M31.2|DMDICD10|LETHAL MIDLINE GRANULOMA|LETALES MITTELLINIENGRANULOM
C2717961|T047|M31.1|DMDICD10|THROMBOTIC MICROANGIOPATHY|THROMBOTISCHE MIKROANGIOPATHIE
C0403529|T047||ICD10CM|HYPERSENSITIVITY ANGIITIS
C2347126|T047||ICD10CM|MICROSCOPIC POLYANGIITIS
C0477585|T047|M31.6|DMDICD10|OTHER GIANT CELL ARTERITIS|SONSTIGE RIESENZELLARTERIITIS
C0343200|T047|M31.5|DMDICD10|GIANT CELL ARTERITIS WITH POLYMYALGIA RHEUMATICA|RIESENZELLARTERIITIS BEI POLYMYALGIA RHEUMATICA
C0039263|T047|M31.4|DMDICD10|AORTIC ARCH SYNDROME [TAKAYASU]|AORTENBOGEN-SYNDROM [TAKAYASU-SYNDROM]
C0477597|T047|M31.9|DMDICD10|NECROTIZING VASCULOPATHY, UNSPECIFIED|NEKROTISIERENDE VASKULOPATHIE, NICHT NAEHER BEZEICHNET
C2895167|T046|M31.8|ICD10CM|OTHER SPECIFIED NECROTIZING VASCULOPATHIES|SEPTIC VASCULITIS
C4270216|T046|T83.031A|ICD10CM|LEAKAGE OF INDWELLING URETHRAL CATHETER, INITIAL ENCOUNTER|LEAKAGE OF INDWELLING URETHRAL CATHETER, INITIAL ENCOUNTER
C4509342|T047|L98.426|ICD10CM|NON-PRESSURE CHRONIC ULCER OF BACK WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULCER OF BACK WITH BONE INVL WITHOUT EVD OF NECR
C2879336|T037|T45.8X2A|ICD10CM|POISONING BY OTHER PRIMARILY SYSTEMIC AND HEMATOLOGICAL AGENTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY OTH PRIM SYS AND HEMATOLOG AGENTS, SLF-HRM, INIT
C3264045|T047|G43.D1|ICD10CM|ABDOMINAL MIGRAINE, INTRACTABLE|ABDOMINAL MIGRAINE, WITH REFRACTORY MIGRAINE
C3264044|T047|G43.D0|ICD10CM|ABDOMINAL MIGRAINE, NOT INTRACTABLE|ABDOMINAL MIGRAINE, NOT INTRACTABLE
C2832178|T037|S06.330A|ICD10CM|CONTUSION AND LACERATION OF CEREBRUM, UNSPECIFIED, WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|CONTUS/LAC CEREB, W/O LOSS OF CONSCIOUSNESS, INIT
C2833375|T037|S12.291A|ICD10CM|OTHER NONDISPLACED FRACTURE OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH NONDISP FX OF THIRD CERVICAL VERTEBRA, INIT FOR CLOS FX
C2833376|T037|S12.291B|ICD10CM|OTHER NONDISPLACED FRACTURE OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH NONDISP FX OF THIRD CERVICAL VERTEBRA, INIT FOR OPN FX
C2891298|T046||ICD10CM|CORNEAL TRANSPLANT INFECTION
C2890682|T037|T84.196A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTERNAL FIXATION DEVICE OF BONE OF RIGHT LOWER LEG, INITIAL ENCOUNTER|MECH COMPL OF INT FIX OF BONE OF RIGHT LOWER LEG, INIT
C2886721|T037|T79.0XXA|ICD10CM|AIR EMBOLISM (TRAUMATIC), INITIAL ENCOUNTER|AIR EMBOLISM (TRAUMATIC), INITIAL ENCOUNTER
C2885207|T037|T61.92XS|ICD10CM|TOXIC EFFECT OF UNSPECIFIED SEAFOOD, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF UNSP SEAFOOD, INTENTIONAL SELF-HARM, SEQUELA
C2884235|T037|T53.2X2A|ICD10CM|TOXIC EFFECT OF TRICHLOROETHYLENE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF TRICHLOROETHYLENE, SELF-HARM, INIT
C2832397|T037|S06.382S|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF BRAINSTEM WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|CONTUS/LAC/HEM BRAINSTEM W LOC OF 31-59 MIN, SEQUELA
C2890076|T037|T82.533A|ICD10CM|LEAKAGE OF BALLOON (COUNTERPULSATION) DEVICE, INITIAL ENCOUNTER|LEAKAGE OF BALLOON (COUNTERPULSATION) DEVICE, INIT ENCNTR
C0477357|T047|G21.8|DMDICD10|OTHER SECONDARY PARKINSONISM|SONSTIGES SEKUNDAERES PARKINSON-SYNDROM
C0030569|T047|G21|DMDICD10|SECONDARY PARKINSONISM, UNSPECIFIED|SEKUNDAERES PARKINSON-SYNDROM
C2884237|T037|T53.2X2S|ICD10CM|TOXIC EFFECT OF TRICHLOROETHYLENE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF TRICHLOROETHYLENE, SELF-HARM, SEQUELA
C0481392|T047|G21.2|DMDICD10|SECONDARY PARKINSONISM DUE TO OTHER EXTERNAL AGENTS|PARKINSON-SYNDROM DURCH SONSTIGE EXOGENE AGENZIEN
C0030568|T047|G21.3|DMDICD10|POSTENCEPHALITIC PARKINSONISM|POSTENZEPHALITISCHES PARKINSON-SYNDROM
C0393568|T047|G21.4|ICD10CM|VASCULAR PARKINSONISM|VASCULAR PARKINSONISM
C4270330|T046|T83.590A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO IMPLANTED URINARY NEUROSTIMULATION DEVICE, INITIAL ENCOUNTER|I/I REACT D/T IMPLANTED URN NSTIM DEV, INITIAL ENCOUNTER
C2887001|T037|T81.532A|ICD10CM|PERFORATION DUE TO FOREIGN BODY ACCIDENTALLY LEFT IN BODY FOLLOWING KIDNEY DIALYSIS, INITIAL ENCOUNTER|PERF DUE TO FB ACC LEFT IN BODY FOL KIDNEY DIALYSIS, INIT
C2889559|T047|M08.23|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, UNSPECIFIED WRIST|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, WRIST
C2887002|T037|T81.532D|ICD10CM|PERFORATION DUE TO FOREIGN BODY ACCIDENTALLY LEFT IN BODY FOLLOWING KIDNEY DIALYSIS, SUBSEQUENT ENCOUNTER|PERF DUE TO FB ACC LEFT IN BODY FOL KIDNEY DIALYSIS, SUBS
C2901220|T046|M84.541A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, RIGHT HAND, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, RIGHT HAND, INIT
C2838409|T037|S32.601B|ICD10CM|UNSPECIFIED FRACTURE OF RIGHT ISCHIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF RIGHT ISCHIUM, INIT FOR OPN FX
C2838408|T037|S32.601A|ICD10CM|UNSPECIFIED FRACTURE OF RIGHT ISCHIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF RIGHT ISCHIUM, INIT FOR CLOS FX
C2887003|T037|T81.532S|ICD10CM|PERFORATION DUE TO FOREIGN BODY ACCIDENTALLY LEFT IN BODY FOLLOWING KIDNEY DIALYSIS, SEQUELA|PERF DUE TO FB ACC LEFT IN BODY FOL KIDNEY DIALYSIS, SEQUELA
C1456308|T048|F31.89|ICD10CM|OTHER BIPOLAR DISORDER|OTHER BIPOLAR DISORDER
C4509114|T048|F31.81|ICD10CM|BIPOLAR II DISORDER|BIPOLAR DISORDER, TYPE 2
C2885815|T037|T63.692A|ICD10CM|TOXIC EFFECT OF CONTACT WITH OTHER VENOMOUS MARINE ANIMALS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFF OF CNTCT W OTH VENOM MARINE ANIMALS, SLF-HRM, INIT
C2876843|T037|T37.2X2A|ICD10CM|POISONING BY ANTIMALARIALS AND DRUGS ACTING ON OTHER BLOOD PROTOZOA, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY ANTIMALARI/DRUGS ACT ON BLD PROTZOA, SLF-HRM, INIT
C2877409|T037|T39.2X2S|ICD10CM|POISONING BY PYRAZOLONE DERIVATIVES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY PYRAZOLONE DERIVATIVES, SELF-HARM, SEQUELA
C2885817|T037|T63.692S|ICD10CM|TOXIC EFFECT OF CONTACT WITH OTHER VENOMOUS MARINE ANIMALS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFF OF CNTCT W OTH VENOM MARINE ANIMALS, SLF-HRM, SQLA
C2876845|T037|T37.2X2S|ICD10CM|POISONING BY ANTIMALARIALS AND DRUGS ACTING ON OTHER BLOOD PROTOZOA, INTENTIONAL SELF-HARM, SEQUELA|POISN BY ANTIMALARI/DRUGS ACT ON BLD PROTZOA, SLF-HRM, SQLA
C4268157|T047|E13.3529|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, UNSPECIFIED EYE|OTH DIAB WITH PROLIF DIAB RTNOP WITH TRCTN DTCH MACULA, UNSP
C2837883|T037|S32.399B|ICD10CM|OTHER FRACTURE OF UNSPECIFIED ILIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTHER FRACTURE OF UNSP ILIUM, INIT ENCNTR FOR OPEN FRACTURE
C2888310|T047|L89.131|ICD10CM|PRESSURE ULCER OF RIGHT LOWER BACK, STAGE 1|PRESSURE ULCER OF RIGHT LOWER BACK, STAGE 1
C2888307|T047||ICD10CM|PRESSURE ULCER OF RIGHT LOWER BACK, UNSTAGEABLE
C2888316|T047|L89.133|ICD10CM|PRESSURE ULCER OF RIGHT LOWER BACK, STAGE 3|PRESSURE ULCER OF RIGHT LOWER BACK, STAGE 3
C2888313|T047|L89.132|ICD10CM|PRESSURE ULCER OF RIGHT LOWER BACK, STAGE 2|PRESSURE ULCER OF RIGHT LOWER BACK, STAGE 2
C4268154|T047|E13.3521|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, RIGHT EYE|OTH DIAB W PROLIF DIAB RTNOP WITH TRCTN DTCH MACULA, R EYE
C4268155|T047|E13.3522|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, LEFT EYE|OTH DIAB W PROLIF DIAB RTNOP WITH TRCTN DTCH MACULA, L EYE
C4268156|T047|E13.3523|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, BILATERAL|OTH DIAB WITH PROLIF DIAB RTNOP WITH TRCTN DTCH MACULA, BI
C2888322|T047|L89.139|ICD10CM|PRESSURE ULCER OF RIGHT LOWER BACK, UNSPECIFIED STAGE|PRESSURE ULCER OF RIGHT LOWER BACK, UNSPECIFIED STAGE
C3161179|T047||ICD10CM|ACQUIRED HEMOPHILIA
C3161181|T047|D68.312|ICD10CM|ANTIPHOSPHOLIPID ANTIBODY WITH HEMORRHAGIC DISORDER|SYSTEMIC LUPUS ERYTHEMATOSUS [SLE] INHIBITOR WITH HEMORRHAGIC DISORDER
C2835182|T037|S22.009A|ICD10CM|UNSPECIFIED FRACTURE OF UNSPECIFIED THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF UNSP THORACIC VERTEBRA, INIT FOR CLOS FX
C2884595|T037|T56.812S|ICD10CM|TOXIC EFFECT OF THALLIUM, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF THALLIUM, INTENTIONAL SELF-HARM, SEQUELA
C2837969|T191|C40.02|ICD10CM|MALIGNANT NEOPLASM OF SCAPULA AND LONG BONES OF LEFT UPPER LIMB|MALIG NEOPLASM OF SCAPULA AND LONG BONES OF LEFT UPPER LIMB
C4270396|T046|T83.721A|ICD10CM|EXPOSURE OF IMPLANTED VAGINAL MESH INTO VAGINA, INITIAL ENCOUNTER|EXPOSURE OF IMPLANTED VAGINAL MESH INTO VAGINA, INIT
C2837967|T191|C40.00|ICD10CM|MALIGNANT NEOPLASM OF SCAPULA AND LONG BONES OF UNSPECIFIED UPPER LIMB|MALIG NEOPLASM OF SCAPULA AND LONG BONES OF UNSP UPPER LIMB
C2837968|T191|C40.01|ICD10CM|MALIGNANT NEOPLASM OF SCAPULA AND LONG BONES OF RIGHT UPPER LIMB|MALIG NEOPLASM OF SCAPULA AND LONG BONES OF RIGHT UPPER LIMB
C2882868|T047|I70.518|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, OTHER EXTREMITY|ATHSCL NONAUT BIO BYPASS OF EXTRM W INTRMT CLAUD, OTH EXTRM
C2882869|T047|I70.519|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, UNSPECIFIED EXTREMITY|ATHSCL NONAUT BIO BYPASS OF EXTRM W INTRMT CLAUD, UNSP EXTRM
C2882865|T047|I70.511|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, RIGHT LEG|ATHSCL NONAUT BIO BYPASS OF EXTRM W INTRMT CLAUD, RIGHT LEG
C2882866|T047|I70.512|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, LEFT LEG|ATHSCL NONAUT BIO BYPASS OF EXTRM W INTRMT CLAUD, LEFT LEG
C2882867|T047|I70.513|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, BILATERAL LEGS|ATHSCL NONAUT BIO BYPASS OF EXTRM W INTRMT CLAUD, BI LEGS
C0003125|T048|F50.00|ICD10CM|ANOREXIA NERVOSA, UNSPECIFIED|ANOREXIA NERVOSA, UNSPECIFIED
C0520608|T048|F50.01|ICD10CM|ANOREXIA NERVOSA, RESTRICTING TYPE|ANOREXIA NERVOSA, RESTRICTING TYPE
C0520609|T048||ICD10CM|ANOREXIA NERVOSA, BINGE EATING/PURGING TYPE
C2876216|T037|T32.77|ICD10CM|CORROSIONS INVOLVING 70-79% OF BODY SURFACE WITH 70-79% THIRD DEGREE CORROSION|CORROS 70-79% OF BODY SURFACE W 70-79% THIRD DEGREE CORROS
C2876215|T037|T32.76|ICD10CM|CORROSIONS INVOLVING 70-79% OF BODY SURFACE WITH 60-69% THIRD DEGREE CORROSION|CORROS 70-79% OF BODY SURFACE W 60-69% THIRD DEGREE CORROS
C2876214|T037|T32.75|ICD10CM|CORROSIONS INVOLVING 70-79% OF BODY SURFACE WITH 50-59% THIRD DEGREE CORROSION|CORROS 70-79% OF BODY SURFACE W 50-59% THIRD DEGREE CORROS
C2876213|T037|T32.74|ICD10CM|CORROSIONS INVOLVING 70-79% OF BODY SURFACE WITH 40-49% THIRD DEGREE CORROSION|CORROS 70-79% OF BODY SURFACE W 40-49% THIRD DEGREE CORROS
C4509322|T047|L97.808|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF UNSPECIFIED LOWER LEG WITH OTHER SPECIFIED SEVERITY|NON-PRS CHRONIC ULCER OTH PRT UNSP LOW LEG WITH OTH SEVERITY
C2888740|T047|L97.809|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF UNSPECIFIED LOWER LEG WITH UNSPECIFIED SEVERITY|NON-PRS CHRONIC ULCER OTH PRT UNSP LOWER LEG W UNSP SEVERITY
C4509321|T047|L97.806|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF UNSPECIFIED LOWER LEG WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OTH PRT UNSP LW LEG W BNE INVL W/O EVD NECR
C2888739|T047|L97.804|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF UNSPECIFIED LOWER LEG WITH NECROSIS OF BONE|NON-PRS CHRONIC ULCER OTH PRT UNSP LOWER LEG W NECROS BONE
C4509320|T047|L97.805|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF UNSPECIFIED LOWER LEG WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OTH PRT UNSP LW LEG W MSL INVL W/O EVD NECR
C2888737|T047|L97.802|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF UNSPECIFIED LOWER LEG WITH FAT LAYER EXPOSED|NON-PRS CHR ULCER OTH PRT UNSP LOW LEG W FAT LAYER EXPOSED
C2888738|T047|L97.803|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF UNSPECIFIED LOWER LEG WITH NECROSIS OF MUSCLE|NON-PRS CHRONIC ULCER OTH PRT UNSP LOWER LEG W NECROS MUSCLE
C2888736|T047|L97.801|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF UNSPECIFIED LOWER LEG LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHR ULCER OTH PRT UNSP LOW LEG LMT TO BRKDWN SKIN
C2883285|T037|T49.0X2S|ICD10CM|POISONING BY LOCAL ANTIFUNGAL, ANTI-INFECTIVE AND ANTI-INFLAMMATORY DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY LOCAL ANTIFUNG/INFECT/INFLAMM DRUGS, SLF-HRM, SQLA
C2883283|T037|T49.0X2A|ICD10CM|POISONING BY LOCAL ANTIFUNGAL, ANTI-INFECTIVE AND ANTI-INFLAMMATORY DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY LOCAL ANTIFUNG/INFECT/INFLAMM DRUGS, SLF-HRM, INIT
C2905760|T037|X78.2XXS|ICD10CM|INTENTIONAL SELF-HARM BY SWORD OR DAGGER, SEQUELA|INTENTIONAL SELF-HARM BY SWORD OR DAGGER, SEQUELA
C2901781|T047|M86.042|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, LEFT HAND|ACUTE HEMATOGENOUS OSTEOMYELITIS, LEFT HAND
C2901780|T047|M86.041|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, RIGHT HAND|ACUTE HEMATOGENOUS OSTEOMYELITIS, RIGHT HAND
C2856949|T037|S72.061B|ICD10CM|DISPLACED ARTICULAR FRACTURE OF HEAD OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPLACED ARTIC FX HEAD OF R FEMUR, INIT FOR OPN FX TYPE I/2
C2856950|T037|S72.061C|ICD10CM|DISPLACED ARTICULAR FRACTURE OF HEAD OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL ARTIC FX HEAD OF R FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2856948|T037|S72.061A|ICD10CM|DISPLACED ARTICULAR FRACTURE OF HEAD OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED ARTICULAR FRACTURE OF HEAD OF RIGHT FEMUR, INIT
C0839932|T047|M86.049|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED HAND|ACUTE HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED HAND
C2834021|T037|S14.148A|ICD10CM|BROWN-SEQUARD SYNDROME AT C8 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|BROWN-SEQUARD SYNDROME AT C8, INIT
C2873876|T047|E05.81|ICD10CM|OTHER THYROTOXICOSIS WITH THYROTOXIC CRISIS OR STORM|OTHER THYROTOXICOSIS WITH THYROTOXIC CRISIS OR STORM
C2873875|T047|E05.80|ICD10CM|OTHER THYROTOXICOSIS WITHOUT THYROTOXIC CRISIS OR STORM|OTHER THYROTOXICOSIS WITHOUT THYROTOXIC CRISIS OR STORM
C4268300|T048|F19.988|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH OTHER PSYCHOACTIVE SUBSTANCE-INDUCED DISORDER|OTHER (OR UNKNOWN) SUBSTANCE-INDUCED OBSESSIVE-COMPULSIVE OR RELATEDDISORDER, WITHOUT USE DISORDER
C4237288|T048|F19.982|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH PSYCHOACTIVE SUBSTANCE-INDUCED SLEEP DISORDER|OTHER (OR UNKNOWN) SUBSTANCE-INDUCED SLEEP DISORDER, WITHOUT USE DISORDER
C4237285|T048|F19.981|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH PSYCHOACTIVE SUBSTANCE-INDUCED SEXUAL DYSFUNCTION|OTHER (OR UNKNOWN) SUBSTANCE-INDUCED SEXUAL DYSFUNCTION, WITHOUT USE DISORDER
C4237264|T048|F19.980|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH PSYCHOACTIVE SUBSTANCE-INDUCED ANXIETY DISORDER|OTHER (OR UNKNOWN) SUBSTANCE-INDUCED ANXIETY DISORDER, WITHOUT USE DISORDER
C2855923|T037|S68.124S|ICD10CM|PARTIAL TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF RIGHT RING FINGER, SEQUELA|PARTIAL TRAUMATIC MCP AMPUTATION OF R RNG FNGR, SEQUELA
C2859152|T037|S73.004A|ICD10CM|UNSPECIFIED DISLOCATION OF RIGHT HIP, INITIAL ENCOUNTER|UNSPECIFIED DISLOCATION OF RIGHT HIP, INITIAL ENCOUNTER
C4268827|T046|M97.01XA|ICD10CM|PERIPROSTHETIC FRACTURE AROUND INTERNAL PROSTHETIC RIGHT HIP JOINT, INITIAL ENCOUNTER|PERIPROSTH FRACTURE AROUND INTERNAL PROSTH R HIP JT, INIT
C0020445|T047|E78.00|ICD10CM|FAMILIAL HYPERCHOLESTEROLEMIA|HYPERBETALIPOPROTEINEMIA
C4270821|T047|E78.00|ICD10CM|PURE HYPERCHOLESTEROLEMIA, UNSPECIFIED|LOW-DENSITY-LIPOPROTEIN-TYPE [LDL] HYPERLIPOPROTEINEMIA
C2874176|T047|E13.65|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH HYPERGLYCEMIA|OTHER SPECIFIED DIABETES MELLITUS WITH HYPERGLYCEMIA
C0348931|T047|E13.69|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATION|OTH DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATION
C2889611|T047|M08.841|ICD10CM|OTHER JUVENILE ARTHRITIS, RIGHT HAND|OTHER JUVENILE ARTHRITIS, RIGHT HAND
C2889612|T047|M08.842|ICD10CM|OTHER JUVENILE ARTHRITIS, LEFT HAND|OTHER JUVENILE ARTHRITIS, LEFT HAND
C3890205|T047|M08.3|DMDICD10|JUVENILE RHEUMATOID POLYARTHRITIS (SERONEGATIVE)|JUVENILE CHRONISCHE ARTHRITIS (SERONEGATIV), POLYARTIKULAER BEGINNENDE FORM
C2882954|T047|I70.648|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF OTHER PART OF LOWER LEG|ATHSCL NONBIOL BYPASS OF LEFT LEG W ULCER OTH PRT LOW LEG
C0409675|T047|M08.1|DMDICD10|JUVENILE ANKYLOSING SPONDYLITIS|JUVENILE SPONDYLITIS ANKYLOSANS
C2874805|T048|F19.182|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE ABUSE WITH PSYCHOACTIVE SUBSTANCE-INDUCED SLEEP DISORDER|OTH PSYCHOACTIVE SUBSTANCE ABUSE W SLEEP DISORDER
C2874804|T048|F19.181|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE ABUSE WITH PSYCHOACTIVE SUBSTANCE-INDUCED SEXUAL DYSFUNCTION|OTH PSYCHOACTIVE SUBSTANCE ABUSE W SEXUAL DYSFUNCTION
C2882955|T047|I70.649|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF UNSPECIFIED SITE|ATHSCL NONBIOL BYPASS OF THE LEFT LEG W ULCER OF UNSP SITE
C2832600|T037|S06.822S|ICD10CM|INJURY OF LEFT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|INJURY OF L INT CAROTID, INTCR W LOC OF 31-59 MIN, SEQUELA
C4316899|T047|E72.04|ICD10CM|CYSTINOSIS|CYSTINOSIS
C0028860|T047||ICD10CM|LOWE'S SYNDROME
C0018609|T047||ICD10CM|HARTNUP'S DISEASE
C0010691|T047|E72.01|ICD10CM|CYSTINURIA|CYSTINURIA
C4268288|T048|F19.188|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE ABUSE WITH OTHER PSYCHOACTIVE SUBSTANCE-INDUCED DISORDER|OTHER (OR UNKNOWN) SUBSTANCE USE DISORDER, MILD, WITH OTHER (OR UNKNOWN) SUBSTANCE INDUCED OBSESSIVE-COMPULSIVE OR RELATED DISORDER
C0010414|T047|B45.9|DMDICD10|CRYPTOCOCCOSIS, UNSPECIFIED|KRYPTOKOKKOSE, NICHT NAEHER BEZEICHNET
C0348251|T047|B45.8|DMDICD10|OTHER FORMS OF CRYPTOCOCCOSIS|SONSTIGE FORMEN DER KRYPTOKOKKOSE
C2838323|T037|S32.483B|ICD10CM|DISPLACED DOME FRACTURE OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISPLACED DOME FRACTURE OF UNSP ACETABULUM, INIT FOR OPN FX
C0276687|T047|B45.7|DMDICD10|DISSEMINATED CRYPTOCOCCOSIS|DISSEMINIERTE KRYPTOKOKKOSE
C2896751|T046|M80.851A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, RIGHT FEMUR, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, RIGHT FEMUR, INIT
C2830239|T047|B45.1|ICD10CM|CEREBRAL CRYPTOCOCCOSIS|CRYPTOCOCCOSIS MENINGOCEREBRALIS
C0276688|T047|B45.0|DMDICD10|PULMONARY CRYPTOCOCCOSIS|KRYPTOKOKKOSE DER LUNGE
C0276690|T047|B45.3|DMDICD10|OSSEOUS CRYPTOCOCCOSIS|KRYPTOKOKKOSE DER KNOCHEN
C0343888|T047|B45.2|DMDICD10|CUTANEOUS CRYPTOCOCCOSIS|KRYPTOKOKKOSE DER HAUT
C2865534|T037|S88.022D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT KNEE LEVEL, LEFT LOWER LEG, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION AT KNEE LEVEL, L LOW LEG, SUBS
C2889364|T047|M05.829|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED ELBOW|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF UNSP ELBOW
C0014804|T047|I73.81|ICD10CM|ERYTHROMELALGIA|ERYTHROMELALGIA
C2901025|T046|M84.461A|ICD10CM|PATHOLOGICAL FRACTURE, RIGHT TIBIA, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, RIGHT TIBIA, INIT ENCNTR FOR FRACTURE
C2889362|T047|M05.821|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT ELBOW|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF RIGHT ELBOW
C2889363|T047|M05.822|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT ELBOW|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF LEFT ELBOW
C2883036|T047|I73.89|ICD10CM|OTHER SPECIFIED PERIPHERAL VASCULAR DISEASES|VASOMOTOR ACROPARESTHESIA [NOTHNAGEL'S TYPE]
C2831434|T037|S02.113S|ICD10CM|UNSPECIFIED OCCIPITAL CONDYLE FRACTURE, SEQUELA|UNSPECIFIED OCCIPITAL CONDYLE FRACTURE, SEQUELA
C2876164|T037|T31.81|ICD10CM|BURNS INVOLVING 80-89% OF BODY SURFACE WITH 10-19% THIRD DEGREE BURNS|BURNS OF 80-89% OF BODY SURFACE W 10-19% THIRD DEGREE BURNS
C2887142|T047|I82.A21|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF RIGHT AXILLARY VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF RIGHT AXILLARY VEIN
C2887143|T047|I82.A22|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF LEFT AXILLARY VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF LEFT AXILLARY VEIN
C2887144|T047|I82.A23|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF AXILLARY VEIN, BILATERAL|CHRONIC EMBOLISM AND THROMBOSIS OF AXILLARY VEIN, BILATERAL
C2876168|T037|T31.85|ICD10CM|BURNS INVOLVING 80-89% OF BODY SURFACE WITH 50-59% THIRD DEGREE BURNS|BURNS OF 80-89% OF BODY SURFACE W 50-59% THIRD DEGREE BURNS
C2876167|T037|T31.84|ICD10CM|BURNS INVOLVING 80-89% OF BODY SURFACE WITH 40-49% THIRD DEGREE BURNS|BURNS OF 80-89% OF BODY SURFACE W 40-49% THIRD DEGREE BURNS
C2876170|T037|T31.87|ICD10CM|BURNS INVOLVING 80-89% OF BODY SURFACE WITH 70-79% THIRD DEGREE BURNS|BURNS OF 80-89% OF BODY SURFACE W 70-79% THIRD DEGREE BURNS
C2887300|T047|I87.311|ICD10CM|CHRONIC VENOUS HYPERTENSION (IDIOPATHIC) WITH ULCER OF RIGHT LOWER EXTREMITY|CHRONIC VENOUS HYPERTENSION W ULCER OF R LOW EXTREM
C2887145|T047|I82.A29|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED AXILLARY VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED AXILLARY VEIN
C2831429|T037|S02.113A|ICD10CM|UNSPECIFIED OCCIPITAL CONDYLE FRACTURE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP OCCIPITAL CONDYLE FRACTURE, INIT FOR CLOS FX
C2882948|T047|I70.642|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF CALF|ATHSCL NONBIOL BYPASS OF THE LEFT LEG W ULCERATION OF CALF
C2831430|T037|S02.113B|ICD10CM|UNSPECIFIED OCCIPITAL CONDYLE FRACTURE, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP OCCIPITAL CONDYLE FRACTURE, INIT FOR OPN FX
C2882949|T047|I70.643|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF ANKLE|ATHSCL NONBIOL BYPASS OF THE LEFT LEG W ULCERATION OF ANKLE
C0477587|T047|M32.8|DMDICD10|OTHER FORMS OF SYSTEMIC LUPUS ERYTHEMATOSUS|SONSTIGE FORMEN DES SYSTEMISCHEN LUPUS ERYTHEMATODES
C2882951|T047|I70.644|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF HEEL AND MIDFOOT|ATHSCL NONBIOL BYPASS OF LEFT LEG W ULCER OF HEEL AND MIDFT
C2902446|T047|M90.562|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, LEFT LOWER LEG|OSTEONECROSIS IN DISEASES CLASSD ELSWHR, LEFT LOWER LEG
C2882953|T047|I70.645|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF OTHER PART OF FOOT|ATHSCL NONBIOL BYPASS OF THE LEFT LEG W ULCER OTH PRT FOOT
C2901531|T046|M84.664A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, LEFT FIBULA, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, LEFT FIBULA, INIT
C0494608|T046|I62.9|DMDICD10|NONTRAUMATIC INTRACRANIAL HEMORRHAGE, UNSPECIFIED|INTRAKRANIELLE BLUTUNG (NICHTTRAUMATISCH), NICHT NAEHER BEZEICHNET
C3263829|T037|S32.82XB|ICD10CM|MULTIPLE FRACTURES OF PELVIS WITHOUT DISRUPTION OF PELVIC RING, INITIAL ENCOUNTER FOR OPEN FRACTURE|MULT FX OF PELVIS W/O DISRUPT OF PELV RING, INIT FOR OPN FX
C2838612|T037|S34.02XS|ICD10CM|CONCUSSION AND EDEMA OF SACRAL SPINAL CORD, SEQUELA|CONCUSSION AND EDEMA OF SACRAL SPINAL CORD, SEQUELA
C2832372|T037|S06.376S|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF CEREBELLUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|CONTUS/LAC/HEM CRBLM W LOC >24 HR W/O RET CONSC W SURV, SQLA
C1318552|T046|I62.1|DMDICD10|NONTRAUMATIC EXTRADURAL HEMORRHAGE|NICHTTRAUMATISCHE EXTRADURALE BLUTUNG
C2901075|T046|M84.473A|ICD10CM|PATHOLOGICAL FRACTURE, UNSPECIFIED ANKLE, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, UNSP ANKLE, INIT ENCNTR FOR FRACTURE
C2838611|T037|S34.02XD|ICD10CM|CONCUSSION AND EDEMA OF SACRAL SPINAL CORD, SUBSEQUENT ENCOUNTER|CONCUSSION AND EDEMA OF SACRAL SPINAL CORD, SUBS ENCNTR
C2838610|T037|S34.02XA|ICD10CM|CONCUSSION AND EDEMA OF SACRAL SPINAL CORD, INITIAL ENCOUNTER|CONCUSSION AND EDEMA OF SACRAL SPINAL CORD, INIT ENCNTR
C0153406|T191|C14.2|DMDICD10|MALIGNANT NEOPLASM OF WALDEYER'S RING|BOESARTIGE NEUBILDUNG: LYMPHATISCHER RACHENRING [WALDEYER]
C4268030|T047|E10.3419|ICD10CM|TYPE 1 DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|TYPE 1 DIAB WITH SEVERE NONP RTNOP WITH MACULAR EDEMA, UNSP
C2901444|T046|M84.639A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, UNSPECIFIED ULNA AND RADIUS, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN OTH DISEASE, UNSP ULNA AND RADIUS, INIT
C4268029|T047|E10.3413|ICD10CM|TYPE 1 DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|TYPE 1 DIAB WITH SEVERE NONP RTNOP WITH MACULAR EDEMA, BI
C4268028|T047|E10.3412|ICD10CM|TYPE 1 DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|TYPE 1 DIAB WITH SEVERE NONP RTNOP WITH MACULAR EDEMA, L EYE
C4268027|T047|E10.3411|ICD10CM|TYPE 1 DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|TYPE 1 DIAB WITH SEVERE NONP RTNOP WITH MACULAR EDEMA, R EYE
C2860215|T037|S79.142A|ICD10CM|SALTER-HARRIS TYPE IV PHYSEAL FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SLTR-HARIS TYPE IV PHYSEAL FX LOWER END OF LEFT FEMUR, INIT
C2896507|T046|M80.021A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, RIGHT HUMERUS, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, R HUMERUS, INIT
C2838386|T037|S32.512A|ICD10CM|FRACTURE OF SUPERIOR RIM OF LEFT PUBIS, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF SUPERIOR RIM OF LEFT PUBIS, INIT FOR CLOS FX
C2869760|T037|S98.012D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT FOOT AT ANKLE LEVEL, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMP OF LEFT FOOT AT ANKLE LEVEL, SUBS
C4270135|T046|T82.828A|ICD10CM|FIBROSIS DUE TO VASCULAR PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|FIBROSIS DUE TO VASCULAR PROSTH DEV/GRFT, INITIAL ENCOUNTER
C2832651|T037|S06.895A|ICD10CM|OTHER SPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, INITIAL ENCOUNTER|INTCRAN INJ W LOC >24 HR W RET CONSC LEV, INIT
C2832653|T037|S06.895S|ICD10CM|OTHER SPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, SEQUELA|INTCRAN INJ W LOC >24 HR W RET CONSC LEV, SEQUELA
C2889488|T047|M06.869|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, UNSPECIFIED KNEE|OTHER SPECIFIED RHEUMATOID ARTHRITIS, UNSPECIFIED KNEE
C2874527|T048|F13.20|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE, UNCOMPLICATED|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE, UNCOMPLICATED
C2874408|T048|F10.92|ICD10CM|ALCOHOL USE, UNSPECIFIED WITH INTOXICATION, UNSPECIFIED|ALCOHOL USE, UNSPECIFIED WITH INTOXICATION
C3263828|T037|S32.82XA|ICD10CM|MULTIPLE FRACTURES OF PELVIS WITHOUT DISRUPTION OF PELVIC RING, INITIAL ENCOUNTER FOR CLOSED FRACTURE|MULTIPLE FX OF PELVIS W/O DISRUPT OF PELVIC RING, INIT
C2874406|T048|F10.920|ICD10CM|ALCOHOL USE, UNSPECIFIED WITH INTOXICATION, UNCOMPLICATED|ALCOHOL USE, UNSPECIFIED WITH INTOXICATION, UNCOMPLICATED
C2874407|T048|F10.921|ICD10CM|ALCOHOL USE, UNSPECIFIED WITH INTOXICATION DELIRIUM|ALCOHOL USE, UNSPECIFIED WITH INTOXICATION DELIRIUM
C2835269|T037|S22.031A|ICD10CM|STABLE BURST FRACTURE OF THIRD THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|STABLE BURST FRACTURE OF THIRD THORACIC VERTEBRA, INIT
C2835270|T037|S22.031B|ICD10CM|STABLE BURST FRACTURE OF THIRD THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|STABLE BURST FX THIRD THOR VERTEBRA, INIT FOR OPN FX
C2837700|T037|S32.120B|ICD10CM|NONDISPLACED ZONE II FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISPLACED ZONE II FRACTURE OF SACRUM, INIT FOR OPN FX
C2837699|T037|S32.120A|ICD10CM|NONDISPLACED ZONE II FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED ZONE II FRACTURE OF SACRUM, INIT FOR CLOS FX
C2832099|T037|S06.311A|ICD10CM|CONTUSION AND LACERATION OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|CONTUS/LAC RIGHT CEREBRUM W LOC OF 30 MINUTES OR LESS, INIT
C2876156|T037|T31.71|ICD10CM|BURNS INVOLVING 70-79% OF BODY SURFACE WITH 10-19% THIRD DEGREE BURNS|BURNS OF 70-79% OF BODY SURFACE W 10-19% THIRD DEGREE BURNS
C2889486|T047|M06.861|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, RIGHT KNEE|OTHER SPECIFIED RHEUMATOID ARTHRITIS, RIGHT KNEE
C0751571|T191|C64-C68|ICD10CM|MALIGNANT NEOPLASM OF URINARY ORGAN, UNSPECIFIED|MALIGNANT NEOPLASMS OF URINARY TRACT (C64-C68)
C2845898|T191|C68.8|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF URINARY ORGANS|PRIMARY MALIGNANT NEOPLASM OF TWO OR MORE CONTIGUOUS SITES OF URINARY ORGANS WHOSE POINT OF ORIGIN CANNOT BE DETERMINED
C2876157|T037|T31.72|ICD10CM|BURNS INVOLVING 70-79% OF BODY SURFACE WITH 20-29% THIRD DEGREE BURNS|BURNS OF 70-79% OF BODY SURFACE W 20-29% THIRD DEGREE BURNS
C2832101|T037|S06.311S|ICD10CM|CONTUSION AND LACERATION OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|CONTUS/LAC R CEREB W LOC OF 30 MINUTES OR LESS, SEQUELA
C0153621|T191|C68.1|DMDICD10|MALIGNANT NEOPLASM OF PARAURETHRAL GLANDS|BOESARTIGE NEUBILDUNG: PARAURETHRALE DRUESE
C0153620|T191|C68.0|DMDICD10|MALIGNANT NEOPLASM OF URETHRA|BOESARTIGE NEUBILDUNG: URETHRA
C4270473|T046|T85.120A|ICD10CM|DISPLACEMENT OF IMPLANTED ELECTRONIC NEUROSTIMULATOR OF BRAIN ELECTRODE (LEAD), INITIAL ENCOUNTER|DISPLACEMENT OF IMPLNT ELEC NSTIM OF BRAIN LEAD, INIT
C2838661|T037|S34.119A|ICD10CM|COMPLETE LESION OF UNSPECIFIED LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION OF UNSP LEVEL OF LUMBAR SPINAL CORD, INIT
C2889487|T047|M06.862|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, LEFT KNEE|OTHER SPECIFIED RHEUMATOID ARTHRITIS, LEFT KNEE
C2838662|T037|S34.119D|ICD10CM|COMPLETE LESION OF UNSPECIFIED LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION OF UNSP LEVEL OF LUMBAR SPINAL CORD, SUBS
C2902374|T047|M89.652|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, LEFT THIGH|OSTEOPATHY AFTER POLIOMYELITIS, LEFT THIGH
C2902373|T047|M89.651|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, RIGHT THIGH|OSTEOPATHY AFTER POLIOMYELITIS, RIGHT THIGH
C2902375|T047|M89.659|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, UNSPECIFIED THIGH|OSTEOPATHY AFTER POLIOMYELITIS, UNSPECIFIED THIGH
C2874505|T048|F12.951|ICD10CM|CANNABIS USE, UNSPECIFIED WITH PSYCHOTIC DISORDER WITH HALLUCINATIONS|CANNABIS USE, UNSP W PSYCHOTIC DISORDER WITH HALLUCINATIONS
C2874504|T048|F12.950|ICD10CM|CANNABIS USE, UNSPECIFIED WITH PSYCHOTIC DISORDER WITH DELUSIONS|CANNABIS USE, UNSP WITH PSYCHOTIC DISORDER WITH DELUSIONS
C2838663|T037|S34.119S|ICD10CM|COMPLETE LESION OF UNSPECIFIED LEVEL OF LUMBAR SPINAL CORD, SEQUELA|COMPLETE LESION OF UNSP LEVEL OF LUMBAR SPINAL CORD, SEQUELA
C4237034|T048|F12.959|ICD10CM|CANNABIS USE, UNSPECIFIED WITH PSYCHOTIC DISORDER, UNSPECIFIED|CANNABIS INDUCED PSYCHOTIC DISORDER, WITHOUT USE DISORDER
C0153570|T191|C53.1|DMDICD10|MALIGNANT NEOPLASM OF EXOCERVIX|BOESARTIGE NEUBILDUNG: EKTOZERVIX
C0153569|T191|C53.0|DMDICD10|MALIGNANT NEOPLASM OF ENDOCERVIX|BOESARTIGE NEUBILDUNG: ENDOZERVIX
C2858268|T037|S72.399A|ICD10CM|OTHER FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF SHAFT OF UNSP FEMUR, INIT FOR CLOS FX
C2858269|T037|S72.399B|ICD10CM|OTHER FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|OTH FX SHAFT OF UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2858270|T037|S72.399C|ICD10CM|OTHER FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|OTH FX SHAFT OF UNSP FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C0007847|T191|C53.9|DMDICD10|MALIGNANT NEOPLASM OF CERVIX UTERI, UNSPECIFIED|BOESARTIGE NEUBILDUNG: CERVIX UTERI, NICHT NAEHER BEZEICHNET
C0348908|T191|C53.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF CERVIX UTERI|BOESARTIGE NEUBILDUNG: CERVIX UTERI, MEHRERE TEILBEREICHE UEBERLAPPEND
C2886000|T037|T65.1X2S|ICD10CM|TOXIC EFFECT OF STRYCHNINE AND ITS SALTS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF STRYCHNINE AND ITS SALTS, SELF-HARM, SEQUELA
C2885984|T037|T65.0X2S|ICD10CM|TOXIC EFFECT OF CYANIDES, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CYANIDES, INTENTIONAL SELF-HARM, SEQUELA
C2885998|T037|T65.1X2A|ICD10CM|TOXIC EFFECT OF STRYCHNINE AND ITS SALTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF STRYCHNINE AND ITS SALTS, SELF-HARM, INIT
C2877359|T037|T39.092S|ICD10CM|POISONING BY SALICYLATES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY SALICYLATES, INTENTIONAL SELF-HARM, SEQUELA
C2885982|T037|T65.0X2A|ICD10CM|TOXIC EFFECT OF CYANIDES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CYANIDES, INTENTIONAL SELF-HARM, INIT ENCNTR
C2890129|T037|T82.6XXA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO CARDIAC VALVE PROSTHESIS, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO CARDIAC VALVE PROSTHESIS, INIT
C2838094|T037|S32.431B|ICD10CM|DISPLACED FRACTURE OF ANTERIOR COLUMN [ILIOPUBIC] OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISP FX OF ANTERIOR COLUMN OF RIGHT ACETAB, INIT FOR OPN FX
C2838093|T037|S32.431A|ICD10CM|DISPLACED FRACTURE OF ANTERIOR COLUMN [ILIOPUBIC] OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF ANTERIOR COLUMN OF RIGHT ACETABULUM, INIT
C2833413|T037|S12.34XB|ICD10CM|TYPE III TRAUMATIC SPONDYLOLISTHESIS OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE III TRAUM SPONDYLOLYSIS OF 4TH CERVCAL VERT, 7THB
C3495801|T047|M31.3|ICD10CM|WEGENER'S GRANULOMATOSIS WITHOUT RENAL INVOLVEMENT|NECROTIZING RESPIRATORY GRANULOMATOSIS
C4268275|T048|F18.14|ICD10CM|INHALANT ABUSE WITH INHALANT-INDUCED MOOD DISORDER|INHALANT USE DISORDER, MILD, WITH INHALANT INDUCED DEPRESSIVE DISORDER
C2842047|T191|C49.21|ICD10CM|MALIGNANT NEOPLASM OF CONNECTIVE AND SOFT TISSUE OF RIGHT LOWER LIMB, INCLUDING HIP|MALIG NEOPLM OF CONN AND SOFT TISS OF R LOW LIMB, INC HIP
C2842046|T191|C49.20|ICD10CM|MALIGNANT NEOPLASM OF CONNECTIVE AND SOFT TISSUE OF UNSPECIFIED LOWER LIMB, INCLUDING HIP|MALIG NEOPLM OF CONN AND SOFT TISS OF UNSP LOW LIMB, INC HIP
C2842048|T191|C49.22|ICD10CM|MALIGNANT NEOPLASM OF CONNECTIVE AND SOFT TISSUE OF LEFT LOWER LIMB, INCLUDING HIP|MALIG NEOPLM OF CONN AND SOFT TISS OF LEFT LOW LIMB, INC HIP
C2887942|T047|K74.69|ICD10CM|OTHER CIRRHOSIS OF LIVER|OTHER CIRRHOSIS OF LIVER
C2853797|T191|C82.12|ICD10CM|FOLLICULAR LYMPHOMA GRADE II, INTRATHORACIC LYMPH NODES|FOLLICULAR LYMPHOMA GRADE II, INTRATHORACIC LYMPH NODES
C2853796|T191|C82.11|ICD10CM|FOLLICULAR LYMPHOMA GRADE II, LYMPH NODES OF HEAD, FACE, AND NECK|FOLLICULAR LYMPHOMA GRADE II, NODES OF HEAD, FACE, AND NECK
C2853795|T191|C82.10|ICD10CM|FOLLICULAR LYMPHOMA GRADE II, UNSPECIFIED SITE|FOLLICULAR LYMPHOMA GRADE II, UNSPECIFIED SITE
C2853802|T191|C82.17|ICD10CM|FOLLICULAR LYMPHOMA GRADE II, SPLEEN|FOLLICULAR LYMPHOMA GRADE II, SPLEEN
C2853801|T191|C82.16|ICD10CM|FOLLICULAR LYMPHOMA GRADE II, INTRAPELVIC LYMPH NODES|FOLLICULAR LYMPHOMA GRADE II, INTRAPELVIC LYMPH NODES
C2853800|T191|C82.15|ICD10CM|FOLLICULAR LYMPHOMA GRADE II, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|FOLICLAR LYMPH GRADE II, NODES OF ING REGION AND LOWER LIMB
C2853799|T191|C82.14|ICD10CM|FOLLICULAR LYMPHOMA GRADE II, LYMPH NODES OF AXILLA AND UPPER LIMB|FOLLICULAR LYMPHOMA GRADE II, NODES OF AXILLA AND UPPER LIMB
C2873882|T047|E08.00|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH HYPEROSMOLARITY WITHOUT NONKETOTIC HYPERGLYCEMIC-HYPEROSMOLAR COMA (NKHHC)|DIAB D/T UNDRL COND W HYPROSM W/O NONKET HYPRGLY-HYPROS COMA
C2873883|T047|E08.01|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH HYPEROSMOLARITY WITH COMA|DIABETES DUE TO UNDERLYING CONDITION W HYPROSM W COMA
C2853804|T191|C82.19|ICD10CM|FOLLICULAR LYMPHOMA GRADE II, EXTRANODAL AND SOLID ORGAN SITES|FOLLICULAR LYMPHOMA GRADE II, EXTRNOD AND SOLID ORGAN SITES
C2853803|T191|C82.18|ICD10CM|FOLLICULAR LYMPHOMA GRADE II, LYMPH NODES OF MULTIPLE SITES|FOLLICULAR LYMPHOMA GRADE II, LYMPH NODES OF MULTIPLE SITES
C0451769|T047|N14.3|DMDICD10|NEPHROPATHY INDUCED BY HEAVY METALS|NEPHROPATHIE DURCH SCHWERMETALLE
C0495053|T046|N14.2|DMDICD10|NEPHROPATHY INDUCED BY UNSPECIFIED DRUG, MEDICAMENT OR BIOLOGICAL SUBSTANCE|NEPHROPATHIE DURCH NICHT NAEHER BEZEICHNETE(S) ARZNEIMITTEL, DROGE ODER BIOLOGISCH AKTIVE SUBSTANZ
C0451767|T046|N14.1|DMDICD10|NEPHROPATHY INDUCED BY OTHER DRUGS, MEDICAMENTS AND BIOLOGICAL SUBSTANCES|NEPHROPATHIE DURCH SONSTIGE ARZNEIMITTEL, DROGEN UND BIOLOGISCH AKTIVE SUBSTANZEN
C0149938|T046|N14.0|DMDICD10|ANALGESIC NEPHROPATHY|ANALGETIKA-NEPHROPATHIE
C0869068|T047|N14.4|DMDICD10|TOXIC NEPHROPATHY, NOT ELSEWHERE CLASSIFIED|TOXISCHE NEPHROPATHIE, ANDERENORTS NICHT KLASSIFIZIERT
C2861605|T191|C92.90|ICD10CM|MYELOID LEUKEMIA, UNSPECIFIED, NOT HAVING ACHIEVED REMISSION|MYELOID LEUKEMIA, UNSPECIFIED, NOT HAVING ACHIEVED REMISSION
C0686593|T191||ICD10AM|MYELOID LEUKEMIA, UNSPECIFIED IN REMISSION
C2349285|T191|C92.92|ICD10CM|MYELOID LEUKEMIA, UNSPECIFIED IN RELAPSE|MYELOID LEUKEMIA, UNSPECIFIED IN RELAPSE
C4269461|T037|S02.620A|ICD10CM|FRACTURE OF SUBCONDYLAR PROCESS OF MANDIBLE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FX SUBCONDYLAR PROCESS OF MANDIBLE, UNSPECIFIED SIDE, INIT
C2888960|T047|M01.X9|ICD10CM|DIRECT INFECTION OF MULTIPLE JOINTS IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIR INFCT OF MULT JOINTS IN INFEC/PARASTC DIS CLASSD ELSWHR
C2888959|T047|M01.X8|ICD10CM|DIRECT INFECTION OF VERTEBRAE IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIRECT INFCT OF VERTEB IN INFEC/PARASTC DIS CLASSD ELSWHR
C2888927|T047|M01.X0|ICD10CM|DIRECT INFECTION OF UNSPECIFIED JOINT IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIR INFCT OF UNSP JOINT IN INFEC/PARASTC DIS CLASSD ELSWHR
C0348932|T047|E13.8|DMDICD10|OTHER SPECIFIED DIABETES MELLITUS WITH UNSPECIFIED COMPLICATIONS|SONSTIGER NAEHER BEZEICHNETER DIABETES MELLITUS: MIT NICHT NAEHER BEZEICHNETEN KOMPLIKATIONEN
C4268380|T047|H35.3213|ICD10CM|EXUDATIVE AGE-RELATED MACULAR DEGENERATION, RIGHT EYE, WITH INACTIVE SCAR|EXUDATIVE AGE-REL MCLR DEGN, RIGHT EYE, WITH INACTIVE SCAR
C4268379|T047|H35.3212|ICD10CM|EXUDATIVE AGE-RELATED MACULAR DEGENERATION, RIGHT EYE, WITH INACTIVE CHOROIDAL NEOVASCULARIZATION|EXDTVE AGE-REL MCLR DEGN, RIGHT EYE, WITH INACT CHRDL NEOVAS
C4268378|T047|H35.3211|ICD10CM|EXUDATIVE AGE-RELATED MACULAR DEGENERATION, RIGHT EYE, WITH ACTIVE CHOROIDAL NEOVASCULARIZATION|EXDTVE AGE-REL MCLR DEGN, RIGHT EYE, WITH ACTV CHRDL NEOVAS
C4268377|T047|H35.3210|ICD10CM|EXUDATIVE AGE-RELATED MACULAR DEGENERATION, RIGHT EYE, STAGE UNSPECIFIED|EXUDATIVE AGE-REL MCLR DEGN, RIGHT EYE, STAGE UNSPECIFIED
C2885043|T037|T60.2X2A|ICD10CM|TOXIC EFFECT OF OTHER INSECTICIDES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF INSECTICIDES, INTENTIONAL SELF-HARM, INIT
C2833234|T037|S12.111A|ICD10CM|POSTERIOR DISPLACED TYPE II DENS FRACTURE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|POSTERIOR DISPLACED TYPE II DENS FRACTURE, INIT FOR CLOS FX
C2833235|T037|S12.111B|ICD10CM|POSTERIOR DISPLACED TYPE II DENS FRACTURE, INITIAL ENCOUNTER FOR OPEN FRACTURE|POSTERIOR DISPLACED TYPE II DENS FRACTURE, INIT FOR OPN FX
C2882108|T047|I21.21|ICD10CM|ST ELEVATION (STEMI) MYOCARDIAL INFARCTION INVOLVING LEFT CIRCUMFLEX CORONARY ARTERY|STEMI INVOLVING LEFT CIRCUMFLEX CORONARY ARTERY
C2885045|T037|T60.2X2S|ICD10CM|TOXIC EFFECT OF OTHER INSECTICIDES, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF INSECTICIDES, INTENTIONAL SELF-HARM, SEQUELA
C2882537|T047|I69.234|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING LEFT NON-DOMINANT SIDE|MONOPLG UPR LMB FOL OTH NTRM INTCRN HEMOR AFF L NONDOM SIDE
C2882536|T047|I69.233|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING RIGHT NON-DOMINANT SIDE|MONOPLG UPR LMB FOL OTH NTRM INTCRN HEMOR AFF R NONDOM SIDE
C2882535|T047|I69.232|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING LEFT DOMINANT SIDE|MONOPLG UPR LMB FOL OTH NTRM INTCRN HEMOR AFF LEFT DOM SIDE
C2882534|T047|I69.231|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING RIGHT DOMINANT SIDE|MONOPLG UPR LMB FOL OTH NTRM INTCRN HEMOR AFF RIGHT DOM SIDE
C2882118|T047|I21.29|ICD10CM|ST ELEVATION (STEMI) MYOCARDIAL INFARCTION INVOLVING OTHER SITES|STEMI INVOLVING OTH SITES
C2882538|T047|I69.239|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING UNSPECIFIED SIDE|MONOPLG UPR LMB FOL OTH NTRM INTCRN HEMOR AFF UNSP SIDE
C2905723|T037|X76.XXXD|ICD10CM|INTENTIONAL SELF-HARM BY SMOKE, FIRE AND FLAMES, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY SMOKE, FIRE AND FLAMES, SUBS ENCNTR
C0477430|T047|G99.2|DMDICD10|MYELOPATHY IN DISEASES CLASSIFIED ELSEWHERE|MYELOPATHIE BEI ANDERENORTS KLASSIFIZIERTEN KRANKHEITEN
C2875409|T047|G99.0|ICD10CM|AUTONOMIC NEUROPATHY IN DISEASES CLASSIFIED ELSEWHERE|AUTONOMIC NEUROPATHY IN DISEASES CLASSIFIED ELSEWHERE
C2905722|T037|X76.XXXA|ICD10CM|INTENTIONAL SELF-HARM BY SMOKE, FIRE AND FLAMES, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY SMOKE, FIRE AND FLAMES, INIT ENCNTR
C2869790|T037|S98.119D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED GREAT TOE, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF UNSP GREAT TOE, SUBS ENCNTR
C3264024|T047|G43.821|ICD10CM|MENSTRUAL MIGRAINE, NOT INTRACTABLE, WITH STATUS MIGRAINOSUS|MENSTRUAL MIGRAINE, NOT INTRACTABLE, WITH STATUS MIGRAINOSUS
C2869791|T037|S98.119S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED GREAT TOE, SEQUELA|COMPLETE TRAUMATIC AMPUTATION OF UNSP GREAT TOE, SEQUELA
C2905724|T037|X76.XXXS|ICD10CM|INTENTIONAL SELF-HARM BY SMOKE, FIRE AND FLAMES, SEQUELA|INTENTIONAL SELF-HARM BY SMOKE, FIRE AND FLAMES, SEQUELA
C2857188|T037|S72.113A|ICD10CM|DISPLACED FRACTURE OF GREATER TROCHANTER OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF GREATER TROCHANTER OF UNSP FEMUR, INIT
C2857189|T037|S72.113B|ICD10CM|DISPLACED FRACTURE OF GREATER TROCHANTER OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF GREATER TROCHANTER OF UNSP FEMR, 7THB
C2857190|T037|S72.113C|ICD10CM|DISPLACED FRACTURE OF GREATER TROCHANTER OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF GREATER TROCHANTER OF UNSP FEMR, 7THC
C2877357|T037|T39.092A|ICD10CM|POISONING BY SALICYLATES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY SALICYLATES, INTENTIONAL SELF-HARM, INIT ENCNTR
C2838629|T037|S34.104D|ICD10CM|UNSPECIFIED INJURY TO L4 LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY TO L4 LEVEL OF LUMBAR SPINAL CORD, SUBS ENCNTR
C2889930|T037|T82.329A|ICD10CM|DISPLACEMENT OF UNSPECIFIED VASCULAR GRAFTS, INITIAL ENCOUNTER|DISPLACEMENT OF UNSPECIFIED VASCULAR GRAFTS, INIT ENCNTR
C2889597|T047|M08.47|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED ANKLE AND FOOT|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, ANKLE AND FOOT
C2878098|T037|T42.2X2S|ICD10CM|POISONING BY SUCCINIMIDES AND OXAZOLIDINEDIONES, INTENTIONAL SELF-HARM, SEQUELA|POISN BY SUCCINIMIDES AND OXAZOLIDINEDIONES, SLF-HRM, SQLA
C2833257|T037|S12.121B|ICD10CM|OTHER NONDISPLACED DENS FRACTURE, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH NONDISPLACED DENS FRACTURE, INIT FOR OPN FX
C2886192|T037|T65.892A|ICD10CM|TOXIC EFFECT OF OTHER SPECIFIED SUBSTANCES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF OTH SUBSTANCES, INTENTIONAL SELF-HARM, INIT
C4270165|T046|T82.856A|ICD10CM|STENOSIS OF PERIPHERAL VASCULAR STENT, INITIAL ENCOUNTER|STENOSIS OF PERIPHERAL VASCULAR STENT, INITIAL ENCOUNTER
C2889595|T047|M08.471|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, RIGHT ANKLE AND FOOT|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, RIGHT ANK/FT
C2889596|T047|M08.472|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, LEFT ANKLE AND FOOT|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, LEFT ANK/FT
C2854118|T191|C91.A2|ICD10CM|MATURE B-CELL LEUKEMIA BURKITT-TYPE, IN RELAPSE|MATURE B-CELL LEUKEMIA BURKITT-TYPE, IN RELAPSE
C2854117|T191|C91.A1|ICD10CM|MATURE B-CELL LEUKEMIA BURKITT-TYPE, IN REMISSION|MATURE B-CELL LEUKEMIA BURKITT-TYPE, IN REMISSION
C2854116|T191|C91.A0|ICD10CM|MATURE B-CELL LEUKEMIA BURKITT-TYPE NOT HAVING ACHIEVED REMISSION|MATURE B-CELL LEUKEMIA BURKITT-TYPE NOT ACHIEVE REMISSION
C2878096|T037|T42.2X2A|ICD10CM|POISONING BY SUCCINIMIDES AND OXAZOLIDINEDIONES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY SUCCINIMIDES AND OXAZOLIDINEDIONES, SELF-HARM, INIT
C0348696|T047|J66.8|DMDICD10|AIRWAY DISEASE DUE TO OTHER SPECIFIC ORGANIC DUSTS|KRANKHEIT DER ATEMWEGE DURCH SONSTIGE NAEHER BEZEICHNETE ORGANISCHE STAEUBE
C2882880|T047|I70.532|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF CALF|ATHSCL NONAUT BIO BYPASS OF THE RIGHT LEG W ULCER OF CALF
C2886194|T037|T65.892S|ICD10CM|TOXIC EFFECT OF OTHER SPECIFIED SUBSTANCES, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF SUBSTANCES, INTENTIONAL SELF-HARM, SEQUELA
C0006866|T047|J66.2|DMDICD10|CANNABINOSIS|CANNABIOSE
C2887471|T047|J66.0|ICD10CM|BYSSINOSIS|AIRWAY DISEASE DUE TO COTTON DUST
C2242894|T047|J66.1|DMDICD10|FLAX-DRESSERS' DISEASE|FLACHSARBEITER-KRANKHEIT
C2883940|T037|T50.Z12S|ICD10CM|POISONING BY IMMUNOGLOBULIN, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY IMMUNOGLOBULIN, INTENTIONAL SELF-HARM, SEQUELA
C2905693|T037|X73.9XXS|ICD10CM|INTENTIONAL SELF-HARM BY UNSPECIFIED LARGER FIREARM DISCHARGE, SEQUELA|SELF-HARM BY UNSP LARGER FIREARM DISCHARGE, SEQUELA
C2887644|T047|K22.719|ICD10CM|BARRETT'S ESOPHAGUS WITH DYSPLASIA, UNSPECIFIED|BARRETT'S ESOPHAGUS WITH DYSPLASIA, UNSPECIFIED
C2835175|T037|S22.008A|ICD10CM|OTHER FRACTURE OF UNSPECIFIED THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF UNSP THORACIC VERTEBRA, INIT FOR CLOS FX
C1334003|T047||ICD10CM|BARRETT'S ESOPHAGUS WITH HIGH GRADE DYSPLASIA
C1334414|T047||ICD10CM|BARRETT'S ESOPHAGUS WITH LOW GRADE DYSPLASIA
C0009447|T047|D83.9|DMDICD10|COMMON VARIABLE IMMUNODEFICIENCY, UNSPECIFIED|VARIABLER IMMUNDEFEKT, NICHT NAEHER BEZEICHNET
C0477327|T047|D83.8|DMDICD10|OTHER COMMON VARIABLE IMMUNODEFICIENCIES|SONSTIGE VARIABLE IMMUNDEFEKTE
C2905692|T037|X73.9XXD|ICD10CM|INTENTIONAL SELF-HARM BY UNSPECIFIED LARGER FIREARM DISCHARGE, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY UNSP LARGER FIREARM DISCHARGE, SUBS
C2905691|T037|X73.9XXA|ICD10CM|INTENTIONAL SELF-HARM BY UNSPECIFIED LARGER FIREARM DISCHARGE, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY UNSP LARGER FIREARM DISCHARGE, INIT
C0451690|T047|D83.1|DMDICD10|COMMON VARIABLE IMMUNODEFICIENCY WITH PREDOMINANT IMMUNOREGULATORY T-CELL DISORDERS|VARIABLER IMMUNDEFEKT MIT UEBERWIEGENDEN IMMUNREGULATORISCHEN T-ZELL-STOERUNGEN
C0451698|T047|D83.0|DMDICD10|COMMON VARIABLE IMMUNODEFICIENCY WITH PREDOMINANT ABNORMALITIES OF B-CELL NUMBERS AND FUNCTION|VARIABLER IMMUNDEFEKT MIT UEBERWIEGENDEN ABWEICHUNGEN DER B-ZELLEN-ZAHL UND -FUNKTION
C0451691|T047|D83.2|DMDICD10|COMMON VARIABLE IMMUNODEFICIENCY WITH AUTOANTIBODIES TO B- OR T-CELLS|VARIABLER IMMUNDEFEKT MIT AUTOANTIKOERPERN GEGEN B- ODER T-ZELLEN
C2890695|T037|T84.210A|ICD10CM|BREAKDOWN (MECHANICAL) OF INTERNAL FIXATION DEVICE OF BONES OF HAND AND FINGERS, INITIAL ENCOUNTER|BREAKDOWN OF INT FIX OF BONES OF HAND AND FINGERS, INIT
C2835824|T037|S24.142S|ICD10CM|BROWN-SEQUARD SYNDROME AT T2-T6 LEVEL OF THORACIC SPINAL CORD, SEQUELA|BROWN-SEQUARD SYNDROME AT T2-T6, SEQUELA
C2856672|T037|S72.026B|ICD10CM|NONDISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF EPIPHY (SEPARATION) (UPPER) OF UNSP FEMR, 7THB
C2856671|T037|S72.026A|ICD10CM|NONDISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF EPIPHY (SEPARATION) (UPPER) OF UNSP FEMR, INIT
C2877995|T037|T41.42XA|ICD10CM|POISONING BY UNSPECIFIED ANESTHETIC, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY UNSP ANESTHETIC, INTENTIONAL SELF-HARM, INIT
C2835823|T037|S24.142D|ICD10CM|BROWN-SEQUARD SYNDROME AT T2-T6 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|BROWN-SEQUARD SYNDROME AT T2-T6, SUBS
C2835822|T037|S24.142A|ICD10CM|BROWN-SEQUARD SYNDROME AT T2-T6 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|BROWN-SEQUARD SYNDROME AT T2-T6, INIT
C2861608|T191|C92.A0|ICD10CM|ACUTE MYELOID LEUKEMIA WITH MULTILINEAGE DYSPLASIA, NOT HAVING ACHIEVED REMISSION|ACUTE MYELOID LEUK W MULTILIN DYSPLASIA, NOT ACHIEVE REMIS
C2861609|T191|C92.A1|ICD10CM|ACUTE MYELOID LEUKEMIA WITH MULTILINEAGE DYSPLASIA, IN REMISSION|ACUTE MYELOID LEUKEMIA W MULTILIN DYSPLASIA, IN REMISSION
C2861610|T191|C92.A2|ICD10CM|ACUTE MYELOID LEUKEMIA WITH MULTILINEAGE DYSPLASIA, IN RELAPSE|ACUTE MYELOID LEUKEMIA W MULTILINEAGE DYSPLASIA, IN RELAPSE
C2887935|T047||ICD10CM|CHRONIC HEPATIC FAILURE WITH COMA
C4268636|T047||ICD10CM|STAGE 1 NECROTIZING ENTEROCOLITIS
C4270811|T047|K55.30|ICD10CM|NECROTIZING ENTEROCOLITIS, UNSPECIFIED|NECROTIZING ENTEROCOLITIS, UNSPECIFIED
C4268638|T047||ICD10CM|STAGE 3 NECROTIZING ENTEROCOLITIS
C4268637|T047||ICD10CM|STAGE 2 NECROTIZING ENTEROCOLITIS
C2858833|T037|S72.456A|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP SUPRCNDL FX W/O INTRCNDL EXTN LOW END UNSP FEMR,INIT
C2858834|T037|S72.456B|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP SUPRCNDL FX W/O INTRCNDL EXTN LOW END UNSP FEMR,7THB
C2858835|T037|S72.456C|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP SUPRCNDL FX W/O INTRCNDL EXTN LOW END UNSP FEMR,7THC
C2838624|T037|S34.103A|ICD10CM|UNSPECIFIED INJURY TO L3 LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY TO L3 LEVEL OF LUMBAR SPINAL CORD, INIT ENCNTR
C2838625|T037|S34.103D|ICD10CM|UNSPECIFIED INJURY TO L3 LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY TO L3 LEVEL OF LUMBAR SPINAL CORD, SUBS ENCNTR
C2889299|T047|M05.619|ICD10CM|RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRIT OF UNSP SHOULDER W INVOLV OF ORGANS AND SYSTEMS
C2838626|T037|S34.103S|ICD10CM|UNSPECIFIED INJURY TO L3 LEVEL OF LUMBAR SPINAL CORD, SEQUELA|UNSP INJURY TO L3 LEVEL OF LUMBAR SPINAL CORD, SEQUELA
C2977645|T033|Z68.43|ICD10CM|BODY MASS INDEX (BMI) 50-59.9 , ADULT|BODY MASS INDEX (BMI) 50-59.9 , ADULT
C2977644|T033|Z68.42|ICD10CM|BODY MASS INDEX (BMI) 45.0-49.9, ADULT|BODY MASS INDEX (BMI) 45.0-49.9, ADULT
C2977647|T033|Z68.45|ICD10CM|BODY MASS INDEX (BMI) 70 OR GREATER, ADULT|BODY MASS INDEX (BMI) 70 OR GREATER, ADULT
C2889298|T047|M05.612|ICD10CM|RHEUMATOID ARTHRITIS OF LEFT SHOULDER WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF L SHOULDER W INVOLV OF ORGANS AND SYSTEMS
C2889297|T047|M05.611|ICD10CM|RHEUMATOID ARTHRITIS OF RIGHT SHOULDER WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF R SHOULDER W INVOLV OF ORGANS AND SYSTEMS
C2977923|T191|C4A.10|ICD10CM|MERKEL CELL CARCINOMA OF UNSPECIFIED EYELID, INCLUDING CANTHUS|MERKEL CELL CARCINOMA OF UNSP EYELID, INCLUDING CANTHUS
C2842051|T191|C4A.11|ICD10CM|MERKEL CELL CARCINOMA OF RIGHT EYELID, INCLUDING CANTHUS|MERKEL CELL CARCINOMA OF RIGHT EYELID, INCLUDING CANTHUS
C2842052|T191|C4A.12|ICD10CM|MERKEL CELL CARCINOMA OF LEFT EYELID, INCLUDING CANTHUS|MERKEL CELL CARCINOMA OF LEFT EYELID, INCLUDING CANTHUS
C2890580|T037|T84.110A|ICD10CM|BREAKDOWN (MECHANICAL) OF INTERNAL FIXATION DEVICE OF RIGHT HUMERUS, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF INT FIX OF RIGHT HUMERUS, INIT
C2832188|T037|S06.332S|ICD10CM|CONTUSION AND LACERATION OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|CONTUS/LAC CEREB, W LOC OF 31-59 MIN, SEQUELA
C2884514|T037|T56.3X2S|ICD10CM|TOXIC EFFECT OF CADMIUM AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CADMIUM AND ITS COMPND, SELF-HARM, SEQUELA
C2832186|T037|S06.332A|ICD10CM|CONTUSION AND LACERATION OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|CONTUS/LAC CEREB, W LOSS OF CONSCIOUSNESS OF 31-59 MIN, INIT
C2884512|T037|T56.3X2A|ICD10CM|TOXIC EFFECT OF CADMIUM AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CADMIUM AND ITS COMPOUNDS, SELF-HARM, INIT
C2875030|T047|G05.4|ICD10CM|MYELITIS IN DISEASES CLASSIFIED ELSEWHERE|MYELITIS IN DISEASES CLASSIFIED ELSEWHERE
C2848415|T037|S58.111A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN ELBOW AND WRIST, RIGHT ARM, INITIAL ENCOUNTER|COMPLETE TRAUM AMP AT LEV BETW ELBOW AND WRIST, R ARM, INIT
C0025306|T047|A39.4|DMDICD10|MENINGOCOCCEMIA, UNSPECIFIED|MENINGOKOKKENSEPSIS, NICHT NAEHER BEZEICHNET
C0343489|T047|A39.3|DMDICD10|CHRONIC MENINGOCOCCEMIA|CHRONISCHE MENINGOKOKKENSEPSIS
C0473877|T047|A39.2|DMDICD10|ACUTE MENINGOCOCCEMIA|AKUTE MENINGOKOKKENSEPSIS
C1403891|T047|A39.1|DMDICD10|WATERHOUSE-FRIDERICHSEN SYNDROME|WATERHOUSE-FRIDERICHSEN-SYNDROM
C2887806|T047|K51.311|ICD10CM|ULCERATIVE (CHRONIC) RECTOSIGMOIDITIS WITH RECTAL BLEEDING|ULCERATIVE (CHRONIC) RECTOSIGMOIDITIS WITH RECTAL BLEEDING
C2874116|T047|E11.622|ICD10CM|TYPE 2 DIABETES MELLITUS WITH OTHER SKIN ULCER|TYPE 2 DIABETES MELLITUS WITH OTHER SKIN ULCER
C2887808|T047|K51.313|ICD10CM|ULCERATIVE (CHRONIC) RECTOSIGMOIDITIS WITH FISTULA|ULCERATIVE (CHRONIC) RECTOSIGMOIDITIS WITH FISTULA
C2887807|T047|K51.312|ICD10CM|ULCERATIVE (CHRONIC) RECTOSIGMOIDITIS WITH INTESTINAL OBSTRUCTION|ULCERATIVE (CHRONIC) RECTOSIGMOIDITIS W INTESTINAL OBST
C2887809|T047|K51.314|ICD10CM|ULCERATIVE (CHRONIC) RECTOSIGMOIDITIS WITH ABSCESS|ULCERATIVE (CHRONIC) RECTOSIGMOIDITIS WITH ABSCESS
C2887811|T047|K51.319|ICD10CM|ULCERATIVE (CHRONIC) RECTOSIGMOIDITIS WITH UNSPECIFIED COMPLICATIONS|ULCERATIVE (CHRONIC) RECTOSIGMOIDITIS W UNSP COMPLICATIONS
C2887810|T047|K51.318|ICD10CM|ULCERATIVE (CHRONIC) RECTOSIGMOIDITIS WITH OTHER COMPLICATION|ULCERATIVE (CHRONIC) RECTOSIGMOIDITIS WITH OTH COMPLICATION
C2874117|T047|E11.628|ICD10CM|TYPE 2 DIABETES MELLITUS WITH OTHER SKIN COMPLICATIONS|TYPE 2 DIABETES MELLITUS WITH OTHER SKIN COMPLICATIONS
C0270733|T047|G23.2|DMDICD10|STRIATONIGRAL DEGENERATION|STRIATONIGRALE DEGENERATION
C0018523|T047|G23.0|DMDICD10|HALLERVORDEN-SPATZ DISEASE|HALLERVORDEN-SPATZ-SYNDROM
C0038868|T047|G23.1|DMDICD10|PROGRESSIVE SUPRANUCLEAR OPHTHALMOPLEGIA [STEELE-RICHARDSON-OLSZEWSKI]|PROGRESSIVE SUPRANUKLEAERE OPHTHALMOPLEGIE [STEELE-RICHARDSON-OLSZEWSKI-SYNDROM]
C2902445|T047|M90.561|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, RIGHT LOWER LEG|OSTEONECROSIS IN DISEASES CLASSD ELSWHR, RIGHT LOWER LEG
C1389280|T046||ICD10CM|OTHER SPECIFIED DEGENERATIVE DISEASES OF BASAL GANGLIA
C0494458|T047|G23.9|DMDICD10|DEGENERATIVE DISEASE OF BASAL GANGLIA, UNSPECIFIED|DEGENERATIVE KRANKHEIT DER BASALGANGLIEN, NICHT NAEHER BEZEICHNET
C2837473|T037|S32.009A|ICD10CM|UNSPECIFIED FRACTURE OF UNSPECIFIED LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF UNSP LUMBAR VERTEBRA, INIT FOR CLOS FX
C2837474|T037|S32.009B|ICD10CM|UNSPECIFIED FRACTURE OF UNSPECIFIED LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF UNSP LUMBAR VERTEBRA, INIT FOR OPN FX
C0837004|T047|E10.36|ICD10AM|TYPE 1 DIABETES MELLITUS WITH DIABETIC CATARACT|TYPE 1 DIABETES MELLITUS WITH DIABETIC CATARACT
C2905815|T037|X83.2XXD|ICD10CM|INTENTIONAL SELF-HARM BY EXPOSURE TO EXTREMES OF COLD, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY EXPOSURE TO EXTREMES OF COLD, SUBS
C0280427|T191|C91.52|ICD10CM|ADULT T-CELL LYMPHOMA/LEUKEMIA (HTLV-1-ASSOCIATED), IN RELAPSE|ADULT T-CELL LYMPHOMA/LEUKEMIA (HTLV-1-ASSOC), IN RELAPSE
C0478099|T046|Q93.5|DMDICD10|OTHER DELETIONS OF PART OF A CHROMOSOME|SONSTIGE DELETIONEN EINES CHROMOSOMENTEILS
C0036221|T191|C96.2|ICD10CM|MAST CELL SARCOMA|MALIGNANT MAST CELL NEOPLASM
C2901292|T046|M84.563A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, RIGHT FIBULA, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, RIGHT FIBULA, INIT
C2905814|T037|X83.2XXA|ICD10CM|INTENTIONAL SELF-HARM BY EXPOSURE TO EXTREMES OF COLD, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY EXPOSURE TO EXTREMES OF COLD, INIT
C2905679|T037|X73.1XXA|ICD10CM|INTENTIONAL SELF-HARM BY HUNTING RIFLE DISCHARGE, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY HUNTING RIFLE DISCHARGE, INIT
C2910109|T019|Q07.03|ICD10CM|ARNOLD-CHIARI SYNDROME WITH SPINA BIFIDA AND HYDROCEPHALUS|ARNOLD-CHIARI SYNDROME WITH SPINA BIFIDA AND HYDROCEPHALUS
C2910108|T019|Q07.02|ICD10CM|ARNOLD-CHIARI SYNDROME WITH HYDROCEPHALUS|ARNOLD-CHIARI SYNDROME WITH HYDROCEPHALUS
C2910107|T019|Q07.01|ICD10CM|ARNOLD-CHIARI SYNDROME WITH SPINA BIFIDA|ARNOLD-CHIARI SYNDROME WITH SPINA BIFIDA
C2910106|T019|Q07.00|ICD10CM|ARNOLD-CHIARI SYNDROME WITHOUT SPINA BIFIDA OR HYDROCEPHALUS|ARNOLD-CHIARI SYNDROME WITHOUT SPINA BIFIDA OR HYDROCEPHALUS
C2833576|T037|S12.591A|ICD10CM|OTHER NONDISPLACED FRACTURE OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH NONDISP FX OF SIXTH CERVICAL VERTEBRA, INIT FOR CLOS FX
C2833577|T037|S12.591B|ICD10CM|OTHER NONDISPLACED FRACTURE OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH NONDISP FX OF SIXTH CERVICAL VERTEBRA, INIT FOR OPN FX
C2895166|T047|M31.31|ICD10CM|WEGENER'S GRANULOMATOSIS WITH RENAL INVOLVEMENT|WEGENER'S GRANULOMATOSIS WITH RENAL INVOLVEMENT
C2857600|T037|S72.23XC|ICD10CM|DISPLACED SUBTROCHANTERIC FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL SUBTROCHNT FX UNSP FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2837973|T191|C40.20|ICD10CM|MALIGNANT NEOPLASM OF LONG BONES OF UNSPECIFIED LOWER LIMB|MALIGNANT NEOPLASM OF LONG BONES OF UNSPECIFIED LOWER LIMB
C2837974|T191|C40.21|ICD10CM|MALIGNANT NEOPLASM OF LONG BONES OF RIGHT LOWER LIMB|MALIGNANT NEOPLASM OF LONG BONES OF RIGHT LOWER LIMB
C2837975|T191|C40.22|ICD10CM|MALIGNANT NEOPLASM OF LONG BONES OF LEFT LOWER LIMB|MALIGNANT NEOPLASM OF LONG BONES OF LEFT LOWER LIMB
C0494723|T047|K25.6|DMDICD10|CHRONIC OR UNSPECIFIED GASTRIC ULCER WITH BOTH HEMORRHAGE AND PERFORATION|ULCUS VENTRICULI: CHRONISCH ODER NICHT NAEHER BEZEICHNET, MIT BLUTUNG UND PERFORATION
C2888287|T047|L89.119|ICD10CM|PRESSURE ULCER OF RIGHT UPPER BACK, UNSPECIFIED STAGE|PRESSURE ULCER OF RIGHT UPPER BACK, UNSPECIFIED STAGE
C0410870|T046|T87.2|DMDICD10|COMPLICATIONS OF OTHER REATTACHED BODY PART|KOMPLIKATIONEN DURCH SONSTIGEN REPLANTIERTEN KOERPERTEIL
C2876194|T037|T32.43|ICD10CM|CORROSIONS INVOLVING 40-49% OF BODY SURFACE WITH 30-39% THIRD DEGREE CORROSION|CORROS 40-49% OF BODY SURFACE W 30-39% THIRD DEGREE CORROS
C2888284|T047|L89.114|ICD10CM|PRESSURE ULCER OF RIGHT UPPER BACK, STAGE 4|PRESSURE ULCER OF RIGHT UPPER BACK, STAGE 4
C2888281|T047|L89.113|ICD10CM|PRESSURE ULCER OF RIGHT UPPER BACK, STAGE 3|PRESSURE ULCER OF RIGHT UPPER BACK, STAGE 3
C2888278|T047|L89.112|ICD10CM|PRESSURE ULCER OF RIGHT UPPER BACK, STAGE 2|PRESSURE ULCER OF RIGHT UPPER BACK, STAGE 2
C2888275|T047|L89.111|ICD10CM|PRESSURE ULCER OF RIGHT UPPER BACK, STAGE 1|PRESSURE ULCER OF RIGHT UPPER BACK, STAGE 1
C2888272|T047||ICD10CM|PRESSURE ULCER OF RIGHT UPPER BACK, UNSTAGEABLE
C2882308|T047|I60.51|ICD10CM|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM RIGHT VERTEBRAL ARTERY|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM R VERTEB ART
C4269511|T037|S02.641B|ICD10CM|FRACTURE OF RAMUS OF RIGHT MANDIBLE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF RAMUS OF RIGHT MANDIBLE, 7THB
C4269510|T037|S02.641A|ICD10CM|FRACTURE OF RAMUS OF RIGHT MANDIBLE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF RAMUS OF RIGHT MANDIBLE, INIT
C2882418|T047|I65.02|ICD10CM|OCCLUSION AND STENOSIS OF LEFT VERTEBRAL ARTERY|OCCLUSION AND STENOSIS OF LEFT VERTEBRAL ARTERY
C4270407|T046|T83.723A|ICD10CM|EXPOSURE OF IMPLANTED URETHRAL BULKING AGENT INTO URETHRA, INITIAL ENCOUNTER|EXPOSURE OF IMPLNT URETHRAL BULKING AGENT INTO URETHRA, INIT
C0476550|T033|Z21|DMDICD10|ASYMPTOMATIC HUMAN IMMUNODEFICIENCY VIRUS [HIV] INFECTION STATUS|ASYMPTOMATISCHE HIV-INFEKTION [HUMANE IMMUNDEFIZIENZ-VIRUSINFEKTION]
C2883734|T037|T50.8X2A|ICD10CM|POISONING BY DIAGNOSTIC AGENTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY DIAGNOSTIC AGENTS, INTENTIONAL SELF-HARM, INIT
C2848443|T037|S58.911S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT FOREARM, LEVEL UNSPECIFIED, SEQUELA|COMPLETE TRAUMATIC AMP OF R FOREARM, LEVEL UNSP, SEQUELA
C2891135|T037|T85.611S|ICD10CM|BREAKDOWN (MECHANICAL) OF INTRAPERITONEAL DIALYSIS CATHETER, SEQUELA|BREAKDOWN OF INTRAPERITONEAL DIALYSIS CATHETER, SEQUELA
C2837919|T037|S32.412A|ICD10CM|DISPLACED FRACTURE OF ANTERIOR WALL OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF ANTERIOR WALL OF LEFT ACETABULUM, INIT
C0271728|T047|E26.1|DMDICD10|SECONDARY HYPERALDOSTERONISM|SEKUNDAERER HYPERALDOSTERONISMUS
C0020428|T047|E26.9|DMDICD10|HYPERALDOSTERONISM, UNSPECIFIED|HYPERALDOSTERONISMUS, NICHT NAEHER BEZEICHNET
C2848441|T037|S58.911A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT FOREARM, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF R FOREARM, LEVEL UNSP, INIT
C0348641|T047|I68.2|DMDICD10|CEREBRAL ARTERITIS IN OTHER DISEASES CLASSIFIED ELSEWHERE|ZEREBRALE ARTERIITIS BEI SONSTIGEN ANDERENORTS KLASSIFIZIERTEN KRANKHEITEN
C2878356|T037|T43.202S|ICD10CM|POISONING BY UNSPECIFIED ANTIDEPRESSANTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY UNSP ANTIDEPRESSANTS, SELF-HARM, SEQUELA
C4509328|T047|L97.828|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF LEFT LOWER LEG WITH OTHER SPECIFIED SEVERITY|NON-PRS CHRONIC ULCER OTH PRT L LOW LEG WITH OTH SEVERITY
C2888752|T047|L97.829|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF LEFT LOWER LEG WITH UNSPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OTH PRT L LOW LEG W UNSP SEVERITY
C2901176|T046|M84.529A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, UNSPECIFIED HUMERUS, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, UNSP HUMERUS, INIT
C2888748|T047|L97.821|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF LEFT LOWER LEG LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHR ULCER OTH PRT L LOW LEG LIMITED TO BRKDWN SKIN
C2888749|T047|L97.822|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF LEFT LOWER LEG WITH FAT LAYER EXPOSED|NON-PRS CHRONIC ULCER OTH PRT L LOW LEG W FAT LAYER EXPOSED
C2888750|T047|L97.823|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF LEFT LOWER LEG WITH NECROSIS OF MUSCLE|NON-PRS CHRONIC ULCER OTH PRT L LOW LEG W NECROSIS OF MUSCLE
C2888751|T047|L97.824|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF LEFT LOWER LEG WITH NECROSIS OF BONE|NON-PRS CHRONIC ULCER OTH PRT L LOW LEG W NECROSIS OF BONE
C4509326|T047|L97.825|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF LEFT LOWER LEG WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OTH PRT L LOW LEG W MSL INVL W/O EVD OF NECR
C4509327|T047|L97.826|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF LEFT LOWER LEG WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OTH PRT L LOW LEG W BNE INVL W/O EVD OF NECR
C2877333|T037|T39.012A|ICD10CM|POISONING BY ASPIRIN, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ASPIRIN, INTENTIONAL SELF-HARM, INIT ENCNTR
C0376329|T047|A81.01|ICD10CM|VARIANT CREUTZFELDT-JAKOB DISEASE|VCJD
C0022336|T047|A81.00|ICD10CM|CREUTZFELDT-JAKOB DISEASE, UNSPECIFIED|CREUTZFELDT-JAKOB DISEASE, UNSPECIFIED
C2900450|T047|A81.09|ICD10CM|OTHER CREUTZFELDT-JAKOB DISEASE|CJD
C2877335|T037|T39.012S|ICD10CM|POISONING BY ASPIRIN, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ASPIRIN, INTENTIONAL SELF-HARM, SEQUELA
C2856759|T037|S72.035B|ICD10CM|NONDISPLACED MIDCERVICAL FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP MIDCERVICAL FX LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C2856758|T037|S72.035A|ICD10CM|NONDISPLACED MIDCERVICAL FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED MIDCERVICAL FRACTURE OF LEFT FEMUR, INIT
C2853798|T191|C82.13|ICD10CM|FOLLICULAR LYMPHOMA GRADE II, INTRA-ABDOMINAL LYMPH NODES|FOLLICULAR LYMPHOMA GRADE II, INTRA-ABDOMINAL LYMPH NODES
C4270435|T046|T83.83XA|ICD10CM|HEMORRHAGE DUE TO GENITOURINARY PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|HEMORRHAGE DUE TO GENITOURINARY PROSTH DEV/GRFT, INIT
C2902101|T046|M87.344|ICD10CM|OTHER SECONDARY OSTEONECROSIS, RIGHT FINGER(S)|OTHER SECONDARY OSTEONECROSIS, RIGHT FINGER(S)
C2885677|T037|T63.452A|ICD10CM|TOXIC EFFECT OF VENOM OF HORNETS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF HORNETS, SELF-HARM, INIT
C2889620|T047|M08.862|ICD10CM|OTHER JUVENILE ARTHRITIS, LEFT KNEE|OTHER JUVENILE ARTHRITIS, LEFT KNEE
C2889619|T047|M08.861|ICD10CM|OTHER JUVENILE ARTHRITIS, RIGHT KNEE|OTHER JUVENILE ARTHRITIS, RIGHT KNEE
C2889621|T047|M08.869|ICD10CM|OTHER JUVENILE ARTHRITIS, UNSPECIFIED KNEE|OTHER JUVENILE ARTHRITIS, UNSPECIFIED KNEE
C2876183|T037|T32.11|ICD10CM|CORROSIONS INVOLVING 10-19% OF BODY SURFACE WITH 10-19% THIRD DEGREE CORROSION|CORROS 10-19% OF BODY SURFACE W 10-19% THIRD DEGREE CORROS
C2874156|T047|E13.49|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH OTHER DIABETIC NEUROLOGICAL COMPLICATION|OTH DIABETES W OTH DIABETIC NEUROLOGICAL COMPLICATION
C2858559|T037|S72.432A|ICD10CM|DISPLACED FRACTURE OF MEDIAL CONDYLE OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF MEDIAL CONDYLE OF LEFT FEMUR, INIT FOR CLOS FX
C2885679|T037|T63.452S|ICD10CM|TOXIC EFFECT OF VENOM OF HORNETS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF HORNETS, SELF-HARM, SEQUELA
C2887939|T047|K74.60|ICD10CM|UNSPECIFIED CIRRHOSIS OF LIVER|UNSPECIFIED CIRRHOSIS OF LIVER
C2874151|T047|E13.40|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC NEUROPATHY, UNSPECIFIED|OTH DIABETES MELLITUS WITH DIABETIC NEUROPATHY, UNSPECIFIED
C0837080|T047|E13.41|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC MONONEUROPATHY|OTH DIABETES MELLITUS WITH DIABETIC MONONEUROPATHY
C2874152|T047|E13.42|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC POLYNEUROPATHY|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC NEURALGIA
C2874154|T047|E13.43|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC AUTONOMIC (POLY)NEUROPATHY|OTH DIABETES MELLITUS W DIABETIC AUTONOMIC (POLY)NEUROPATHY
C2874155|T047|E13.44|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC AMYOTROPHY|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC AMYOTROPHY
C2889370|T047|M05.842|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HAND|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HAND
C2889369|T047|M05.841|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT HAND|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF RIGHT HAND
C2832014|T037|S06.2X0S|ICD10CM|DIFFUSE TRAUMATIC BRAIN INJURY WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|DIFFUSE TBI W/O LOSS OF CONSCIOUSNESS, SEQUELA
C2889371|T047|M05.84|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED HAND|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF HAND
C4268071|T047|E11.3219|ICD10CM|TYPE 2 DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|TYPE 2 DIAB WITH MILD NONP RTNOP WITH MACULAR EDEMA, UNSP
C0270788|T047|G83.9|DMDICD10|PARALYTIC SYNDROME, UNSPECIFIED|LAEHMUNGSSYNDROM, NICHT NAEHER BEZEICHNET
C0694548|T047|J45.991|ICD10CM|COUGH VARIANT ASTHMA|COUGH VARIANT ASTHMA
C0015263|T047||ICD10CM|EXERCISE INDUCED BRONCHOSPASM
C0154701|T047|G83.0|DMDICD10|DIPLEGIA OF UPPER LIMBS|DIPLEGIE DER OBEREN EXTREMITAETEN
C2833863|T037|S14.105D|ICD10CM|UNSPECIFIED INJURY AT C5 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY AT C5 LEVEL OF CERVICAL SPINAL CORD, SUBS ENCNTR
C2875357|T046|G83.4|ICD10CM|CAUDA EQUINA SYNDROME|NEUROGENIC BLADDER DUE TO CAUDA EQUINA SYNDROME
C2887466|T047|J45.998|ICD10CM|OTHER ASTHMA|OTHER ASTHMA
C2833862|T037|S14.105A|ICD10CM|UNSPECIFIED INJURY AT C5 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY AT C5 LEVEL OF CERVICAL SPINAL CORD, INIT ENCNTR
C4087263|T048|F34.1|ICD10CM|DYSTHYMIC DISORDER|PERSISTENT DEPRESSIVE DISORDER
C0010598|T048|F34.0|DMDICD10|CYCLOTHYMIC DISORDER|ZYKLOTHYMIA
C0349224|T048|F34|DMDICD10|PERSISTENT MOOD [AFFECTIVE] DISORDER, UNSPECIFIED|ANHALTENDE AFFEKTIVE STOERUNGEN
C2833864|T037|S14.105S|ICD10CM|UNSPECIFIED INJURY AT C5 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|UNSP INJURY AT C5 LEVEL OF CERVICAL SPINAL CORD, SEQUELA
C2882297|T046|I60.2|ICD10CM|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM ANTERIOR COMMUNICATING ARTERY|NTRM SUBARACH HEMORRHAGE FROM ANTERIOR COMMUNICATING ARTERY
C2882305|T047|I60.4|ICD10CM|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM BASILAR ARTERY|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM BASILAR ARTERY
C2875171|T047|G43.619|ICD10CM|PERSISTENT MIGRAINE AURA WITH CEREBRAL INFARCTION, INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|PERST MIGRAINE AURA W CEREBRAL INFRC, NTRCT, W/O STAT MIGR
C2882310|T047|I60.6|ICD10CM|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM OTHER INTRACRANIAL ARTERIES|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM OTH INTRACRAN ART
C1410400|T047|I60.9|ICD10CM|NONTRAUMATIC SUBARACHNOID HEMORRHAGE, UNSPECIFIED|NONTRAUMATIC SUBARACHNOID HEMORRHAGE, UNSPECIFIED
C2882316|T047|I60.8|ICD10CM|OTHER NONTRAUMATIC SUBARACHNOID HEMORRHAGE|OTHER NONTRAUMATIC SUBARACHNOID HEMORRHAGE
C2875170|T047|G43.611|ICD10CM|PERSISTENT MIGRAINE AURA WITH CEREBRAL INFARCTION, INTRACTABLE, WITH STATUS MIGRAINOSUS|PERST MIGRAINE AURA W CEREBRAL INFRC, NTRCT, W STAT MIGR
C2833308|T037|S12.191A|ICD10CM|OTHER NONDISPLACED FRACTURE OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH NONDISP FX OF SECOND CERVICAL VERTEBRA, INIT FOR CLOS FX
C2833309|T037|S12.191B|ICD10CM|OTHER NONDISPLACED FRACTURE OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH NONDISP FX OF SECOND CERVICAL VERTEBRA, INIT FOR OPN FX
C0268247|T047||ICD10CM|NIEMANN-PICK DISEASE TYPE D
C0220756|T047||ICD10CM|NIEMANN-PICK DISEASE TYPE C
C0268243|T047||ICD10CM|NIEMANN-PICK DISEASE TYPE B
C0268242|T047||ICD10CM|NIEMANN-PICK DISEASE TYPE A
C0028064|T047|E75.249|ICD10CM|NIEMANN-PICK DISEASE, UNSPECIFIED|NIEMANN-PICK DISEASE, UNSPECIFIED
C2874273|T047|E75.248|ICD10CM|OTHER NIEMANN-PICK DISEASE|OTHER NIEMANN-PICK DISEASE
C2832513|T037|S06.6X1A|ICD10CM|TRAUMATIC SUBARACHNOID HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|TRAUM SUBRAC HEM W LOC OF 30 MINUTES OR LESS, INIT
C2901061|T046|M84.471A|ICD10CM|PATHOLOGICAL FRACTURE, RIGHT ANKLE, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, RIGHT ANKLE, INIT ENCNTR FOR FRACTURE
C2882681|T046|I69.969|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING UNSPECIFIED SIDE|OTH PARLYT SYNDROME FOL UNSP CEREBVASC DISEASE AFF UNSP SIDE
C4270439|T046|T83.84XA|ICD10CM|PAIN DUE TO GENITOURINARY PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|PAIN DUE TO GENITOURINARY PROSTH DEV/GRFT, INITIAL ENCOUNTER
C0840138|T047|M89.69|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, MULTIPLE SITES|OSTEOPATHY AFTER POLIOMYELITIS, MULTIPLE SITES
C2889188|T047|M05.262|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT KNEE|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889187|T047|M05.261|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT KNEE|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889189|T047|M05.269|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSP KNEE
C0348806|T047|J85.1|DMDICD10|ABSCESS OF LUNG WITH PNEUMONIA|ABSZESS DER LUNGE MIT PNEUMONIE
C0494682|T047|J85.0|DMDICD10|GANGRENE AND NECROSIS OF LUNG|GANGRAEN UND NEKROSE DER LUNGE
C0155909|T047|J85.3|DMDICD10|ABSCESS OF MEDIASTINUM|ABSZESS DES MEDIASTINUMS
C0494683|T047|J85.2|DMDICD10|ABSCESS OF LUNG WITHOUT PNEUMONIA|ABSZESS DER LUNGE OHNE PNEUMONIE
C2887492|T046|J95.01|ICD10CM|HEMORRHAGE FROM TRACHEOSTOMY STOMA|HEMORRHAGE FROM TRACHEOSTOMY STOMA
C0155921|T046|J95.00|ICD10CM|UNSPECIFIED TRACHEOSTOMY COMPLICATION|UNSPECIFIED TRACHEOSTOMY COMPLICATION
C2887495|T046|J95.03|ICD10CM|MALFUNCTION OF TRACHEOSTOMY STOMA|MALFUNCTION OF TRACHEOSTOMY STOMA
C2711621|T047|J95.02|ICD10CM|INFECTION OF TRACHEOSTOMY STOMA|INFECTION OF TRACHEOSTOMY STOMA
C0695238|T046|J95.09|ICD10CM|OTHER TRACHEOSTOMY COMPLICATION|OTHER TRACHEOSTOMY COMPLICATION
C4269462|T037|S02.620B|ICD10CM|FRACTURE OF SUBCONDYLAR PROCESS OF MANDIBLE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FX SUBCONDYLAR PROCESS OF MANDIBLE, UNSPECIFIED SIDE, 7THB
C2845976|T191|C7A.00|ICD10CM|MALIGNANT CARCINOID TUMOR OF UNSPECIFIED SITE|MALIGNANT CARCINOID TUMOR OF UNSPECIFIED SITE
C2886349|T037|T71.122S|ICD10CM|ASPHYXIATION DUE TO PLASTIC BAG, INTENTIONAL SELF-HARM, SEQUELA|ASPHYXIATION DUE TO PLASTIC BAG, SELF-HARM, SEQUELA
C2885933|T037|T63.92XA|ICD10CM|TOXIC EFFECT OF CONTACT WITH UNSPECIFIED VENOMOUS ANIMAL, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CONTACT W UNSP VENOM ANIMAL, SLF-HRM, INIT
C4268795|T046|M84.757A|ICD10CM|COMPLETE OBLIQUE ATYPICAL FEMORAL FRACTURE, RIGHT LEG, INITIAL ENCOUNTER FOR FRACTURE|COMPLETE OBLIQUE ATYPICAL FEMORAL FRACTURE, RIGHT LEG, INIT
C2876169|T037|T31.86|ICD10CM|BURNS INVOLVING 80-89% OF BODY SURFACE WITH 60-69% THIRD DEGREE BURNS|BURNS OF 80-89% OF BODY SURFACE W 60-69% THIRD DEGREE BURNS
C2860012|T037|S78.121S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN RIGHT HIP AND KNEE, SEQUELA|PARTIAL TRAUMATIC AMP AT LEVEL BETW R HIP AND KNEE, SEQUELA
C2885935|T037|T63.92XS|ICD10CM|TOXIC EFFECT OF CONTACT WITH UNSPECIFIED VENOMOUS ANIMAL, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CNTCT W UNSP VENOM ANIMAL, SLF-HRM, SEQUELA
C2855893|T037|S68.117S|ICD10CM|COMPLETE TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF LEFT LITTLE FINGER, SEQUELA|COMPLETE TRAUMATIC MCP AMP OF L LITTLE FINGER, SEQUELA
C2891223|T037|T85.71XA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO PERITONEAL DIALYSIS CATHETER, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO PERITON DIALYSIS CATHETER, INIT
C2891224|T037|T85.71XD|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO PERITONEAL DIALYSIS CATHETER, SUBSEQUENT ENCOUNTER|INFECT/INFLM REACTION DUE TO PERITON DIALYSIS CATHETER, SUBS
C2837467|T037|S32.008B|ICD10CM|OTHER FRACTURE OF UNSPECIFIED LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF UNSP LUMBAR VERTEBRA, INIT FOR OPN FX
C2901270|T046|M84.559A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, HIP, UNSPECIFIED, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, HIP, UNSP, INIT
C2878871|T037|T44.5X2S|ICD10CM|POISONING BY PREDOMINANTLY BETA-ADRENORECEPTOR AGONISTS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY PREDOM BETA-ADRENOCPT AGONISTS, SELF-HARM, SEQUELA
C2891225|T037|T85.71XS|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO PERITONEAL DIALYSIS CATHETER, SEQUELA|INFECT/INFLM REACTION DUE TO PERITON DIALYSIS CATH, SEQUELA
C2878869|T037|T44.5X2A|ICD10CM|POISONING BY PREDOMINANTLY BETA-ADRENORECEPTOR AGONISTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY PREDOM BETA-ADRENOCPT AGONISTS, SELF-HARM, INIT
C2902366|T047|M89.631|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, RIGHT FOREARM|OSTEOPATHY AFTER POLIOMYELITIS, RIGHT FOREARM
C2902367|T047|M89.632|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, LEFT FOREARM|OSTEOPATHY AFTER POLIOMYELITIS, LEFT FOREARM
C2876171|T037|T31.88|ICD10CM|BURNS INVOLVING 80-89% OF BODY SURFACE WITH 80-89% THIRD DEGREE BURNS|BURNS OF 80-89% OF BODY SURFACE W 80-89% THIRD DEGREE BURNS
C2902368|T047|M89.639|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, UNSPECIFIED FOREARM|OSTEOPATHY AFTER POLIOMYELITIS, UNSPECIFIED FOREARM
C0840146|T047|M89.68|ICD10AM|OSTEOPATHY AFTER POLIOMYELITIS, OTHER SITE|OSTEOPATHY AFTER POLIOMYELITIS, OTHER SITE
C4269466|T037|S02.620S|ICD10CM|FRACTURE OF SUBCONDYLAR PROCESS OF MANDIBLE, UNSPECIFIED SIDE, SEQUELA|FX SUBCONDYLAR PROCESS OF MANDIBLE, UNSP SIDE, SEQUELA
C2905784|T037|X81.1XXS|ICD10CM|INTENTIONAL SELF-HARM BY JUMPING OR LYING IN FRONT OF (SUBWAY) TRAIN, SEQUELA|SLF-HRM BY JUMPING OR LYING IN FRONT OF TRAIN, SEQUELA
C0040128|T047|E07.9|DMDICD10|DISORDER OF THYROID, UNSPECIFIED|KRANKHEIT DER SCHILDDRUESE, NICHT NAEHER BEZEICHNET
C2901306|T046|M84.569A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, UNSPECIFIED TIBIA AND FIBULA, INITIAL ENCOUNTER FOR FRACTURE|PATH FX IN NEOPLTC DISEASE, UNSP TIBIA AND FIBULA, INIT
C0342190|T047|E07.0|ICD10CM|HYPERSECRETION OF CALCITONIN|C-CELL HYPERPLASIA OF THYROID
C2873879|T047|E07.1|ICD10CM|DYSHORMOGENETIC GOITER|FAMILIAL DYSHORMOGENETIC GOITER
C2905782|T037|X81.1XXA|ICD10CM|INTENTIONAL SELF-HARM BY JUMPING OR LYING IN FRONT OF (SUBWAY) TRAIN, INITIAL ENCOUNTER|SLF-HRM BY JUMPING OR LYING IN FRONT OF (SUBWAY) TRAIN, INIT
C2905783|T037|X81.1XXD|ICD10CM|INTENTIONAL SELF-HARM BY JUMPING OR LYING IN FRONT OF (SUBWAY) TRAIN, SUBSEQUENT ENCOUNTER|SLF-HRM BY JUMPING OR LYING IN FRONT OF (SUBWAY) TRAIN, SUBS
C1399358|T047||ICD10CM|PARKINSON'S DISEASE
C2838107|T037|S32.433A|ICD10CM|DISPLACED FRACTURE OF ANTERIOR COLUMN [ILIOPUBIC] OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF ANTERIOR COLUMN OF UNSP ACETABULUM, INIT
C2838108|T037|S32.433B|ICD10CM|DISPLACED FRACTURE OF ANTERIOR COLUMN [ILIOPUBIC] OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISP FX OF ANTERIOR COLUMN OF UNSP ACETAB, INIT FOR OPN FX
C2845966|T191|C79.02|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF LEFT KIDNEY AND RENAL PELVIS|SECONDARY MALIGNANT NEOPLASM OF LEFT KIDNEY AND RENAL PELVIS
C2845964|T191|C79.00|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF UNSPECIFIED KIDNEY AND RENAL PELVIS|SECONDARY MALIGNANT NEOPLASM OF UNSP KIDNEY AND RENAL PELVIS
C2845965|T191|C79.01|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF RIGHT KIDNEY AND RENAL PELVIS|SECONDARY MALIGNANT NEOPLASM OF R KIDNEY AND RENAL PELVIS
C2878561|T037|T43.602A|ICD10CM|POISONING BY UNSPECIFIED PSYCHOSTIMULANTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY UNSP PSYCHOSTIMULANTS, SELF-HARM, INIT
C2861645|T191|C95.00|ICD10CM|ACUTE LEUKEMIA OF UNSPECIFIED CELL TYPE NOT HAVING ACHIEVED REMISSION|ACUTE LEUKEMIA OF UNSP CELL TYPE NOT ACHIEVE REMISSION
C0686586|T191||ICD10AM|ACUTE LEUKEMIA OF UNSPECIFIED CELL TYPE, IN REMISSION
C2349305|T191|C95.02|ICD10CM|ACUTE LEUKEMIA OF UNSPECIFIED CELL TYPE, IN RELAPSE|ACUTE LEUKEMIA OF UNSPECIFIED CELL TYPE, IN RELAPSE
C2890716|T037|T84.223A|ICD10CM|DISPLACEMENT OF INTERNAL FIXATION DEVICE OF BONES OF FOOT AND TOES, INITIAL ENCOUNTER|DISPLACEMENT OF INT FIX OF BONES OF FOOT AND TOES, INIT
C2878563|T037|T43.602S|ICD10CM|POISONING BY UNSPECIFIED PSYCHOSTIMULANTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY UNSP PSYCHOSTIMULANTS, SELF-HARM, SEQUELA
C2883558|T037|T50.1X2A|ICD10CM|POISONING BY LOOP [HIGH-CEILING] DIURETICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY LOOP DIURETICS, INTENTIONAL SELF-HARM, INIT
C2890630|T037|T84.123A|ICD10CM|DISPLACEMENT OF INTERNAL FIXATION DEVICE OF BONE OF LEFT FOREARM, INITIAL ENCOUNTER|DISPLACEMENT OF INT FIX OF BONE OF LEFT FOREARM, INIT
C4237393|T048|F13.980|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED ANXIETY DISORDER|SEDATIVE, HYPNOTIC, OR ANXIOLYTIC-INDUCED ANXIETY DISORDER, WITHOUT USE DISORDER
C4237413|T048|F13.982|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED SLEEP DISORDER|SEDATIVE, HYPNOTIC, OR ANXIOLYTIC-INDUCED SLEEP DISORDER, WITHOUT USE DISORDER
C2853710|T191|C80.1|ICD10CM|MALIGNANT (PRIMARY) NEOPLASM, UNSPECIFIED|MALIGNANT (PRIMARY) NEOPLASM, UNSPECIFIED
C2845988|T191|C80.0|ICD10CM|DISSEMINATED MALIGNANT NEOPLASM, UNSPECIFIED|DISSEMINATED MALIGNANT NEOPLASM, UNSPECIFIED
C2349259|T191||ICD10CM|MALIGNANT NEOPLASM ASSOCIATED WITH TRANSPLANTED ORGAN
C2896640|T046|M80.08XA|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, VERTEBRA(E), INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, VERTEBRA(E), INIT
C2831458|T037|S02.19XS|ICD10CM|OTHER FRACTURE OF BASE OF SKULL, SEQUELA|OTHER FRACTURE OF BASE OF SKULL, SEQUELA
C2901285|T046|M84.562A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, LEFT TIBIA, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, LEFT TIBIA, INIT
C2901430|T047|M84.633A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, RIGHT RADIUS, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, RIGHT RADIUS, INIT
C2865565|T037|S88.129S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, UNSPECIFIED LOWER LEG, SEQUELA|PART TRAUM AMP AT LEV BETW KNEE AND ANKL, UNSP LOW LEG, SQLA
C2858458|T037|S72.422B|ICD10CM|DISPLACED FRACTURE OF LATERAL CONDYLE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF LATERAL CONDYLE OF L FEMR, 7THB
C4268387|T047|H35.3231|ICD10CM|EXUDATIVE AGE-RELATED MACULAR DEGENERATION, BILATERAL, WITH ACTIVE CHOROIDAL NEOVASCULARIZATION|EXUDATIVE AGE-REL MCLR DEGN, BI, WITH ACTV CHRDL NEOVAS
C4268386|T047|H35.3230|ICD10CM|EXUDATIVE AGE-RELATED MACULAR DEGENERATION, BILATERAL, STAGE UNSPECIFIED|EXUDATIVE AGE-REL MCLR DEGN, BILATERAL, STAGE UNSPECIFIED
C4268389|T047|H35.3233|ICD10CM|EXUDATIVE AGE-RELATED MACULAR DEGENERATION, BILATERAL, WITH INACTIVE SCAR|EXUDATIVE AGE-REL MCLR DEGN, BILATERAL, WITH INACTIVE SCAR
C4268388|T047|H35.3232|ICD10CM|EXUDATIVE AGE-RELATED MACULAR DEGENERATION, BILATERAL, WITH INACTIVE CHOROIDAL NEOVASCULARIZATION|EXUDATIVE AGE-REL MCLR DEGN, BI, WITH INACT CHRDL NEOVAS
C2882546|T047|I69.251|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING RIGHT DOMINANT SIDE|HEMIPLGA FOL OTH NTRM INTCRN HEMOR AFF RIGHT DOMINANT SIDE
C2882548|T047|I69.253|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING RIGHT NON-DOMINANT SIDE|HEMIPLGA FOL OTH NTRM INTCRN HEMOR AFF RIGHT NONDOM SIDE
C2882547|T047|I69.252|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING LEFT DOMINANT SIDE|HEMIPLGA FOL OTH NTRM INTCRN HEMOR AFF LEFT DOMINANT SIDE
C2882549|T047|I69.254|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING LEFT NON-DOMINANT SIDE|HEMIPLGA FOL OTH NTRM INTCRN HEMOR AFF LEFT NONDOM SIDE
C2882098|T047|I21.09|ICD10CM|ST ELEVATION (STEMI) MYOCARDIAL INFARCTION INVOLVING OTHER CORONARY ARTERY OF ANTERIOR WALL|STEMI INVOLVING OTH CORONARY ARTERY OF ANTERIOR WALL
C2882550|T047|I69.259|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING UNSPECIFIED SIDE|HEMIPLGA FOLLOWING OTH NTRM INTCRN HEMOR AFFECTING UNSP SIDE
C2882093|T047|I21.02|ICD10CM|ST ELEVATION (STEMI) MYOCARDIAL INFARCTION INVOLVING LEFT ANTERIOR DESCENDING CORONARY ARTERY|STEMI INVOLVING LEFT ANTERIOR DESCENDING CORONARY ARTERY
C2882091|T047|I21.01|ICD10CM|ST ELEVATION (STEMI) MYOCARDIAL INFARCTION INVOLVING LEFT MAIN CORONARY ARTERY|STEMI INVOLVING LEFT MAIN CORONARY ARTERY
C2835761|T037|S24.102D|ICD10CM|UNSPECIFIED INJURY AT T2-T6 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY AT T2-T6 LEVEL OF THORACIC SPINAL CORD, SUBS
C2856094|T037|S68.719A|ICD10CM|COMPLETE TRAUMATIC TRANSMETACARPAL AMPUTATION OF UNSPECIFIED HAND, INITIAL ENCOUNTER|COMPLETE TRAUMATIC TRANSMETCRPL AMP OF UNSP HAND, INIT
C2832505|T037|S06.5X9A|ICD10CM|TRAUMATIC SUBDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|TRAUM SUBDR HEM W LOC OF UNSP DURATION, INIT
C4268135|T047|E13.3313|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|OTH DIABETES WITH MODERATE NONP RTNOP WITH MACULAR EDEMA, BI
C4268134|T047|E13.3312|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|OTH DIAB WITH MODERATE NONP RTNOP WITH MACULAR EDEMA, L EYE
C4268133|T047|E13.3311|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|OTH DIAB WITH MODERATE NONP RTNOP WITH MACULAR EDEMA, R EYE
C4268136|T047|E13.3319|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|OTH DIAB WITH MODERATE NONP RTNOP WITH MACULAR EDEMA, UNSP
C2856096|T037|S68.719S|ICD10CM|COMPLETE TRAUMATIC TRANSMETACARPAL AMPUTATION OF UNSPECIFIED HAND, SEQUELA|COMPLETE TRAUMATIC TRANSMETCRPL AMP OF UNSP HAND, SEQUELA
C2888835|T047|M00.129|ICD10CM|PNEUMOCOCCAL ARTHRITIS, UNSPECIFIED ELBOW|PNEUMOCOCCAL ARTHRITIS, UNSPECIFIED ELBOW
C2888834|T047|M00.122|ICD10CM|PNEUMOCOCCAL ARTHRITIS, LEFT ELBOW|PNEUMOCOCCAL ARTHRITIS, LEFT ELBOW
C2888833|T047|M00.121|ICD10CM|PNEUMOCOCCAL ARTHRITIS, RIGHT ELBOW|PNEUMOCOCCAL ARTHRITIS, RIGHT ELBOW
C4268122|T047|E11.37X2|ICD10CM|TYPE 2 DIABETES MELLITUS WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, LEFT EYE|TYPE 2 DIAB WITH DIAB MCLR EDEMA, RESOLVED FOL TRTMT, L EYE
C4268123|T047|E11.37X3|ICD10CM|TYPE 2 DIABETES MELLITUS WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, BILATERAL|TYPE 2 DIAB WITH DIAB MACULAR EDEMA, RESOLVED FOL TRTMT, BI
C4268121|T047|E11.37X1|ICD10CM|TYPE 2 DIABETES MELLITUS WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, RIGHT EYE|TYPE 2 DIAB WITH DIAB MCLR EDEMA, RESOLVED FOL TRTMT, R EYE
C4268124|T047|E11.37X9|ICD10CM|TYPE 2 DIABETES MELLITUS WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, UNSPECIFIED EYE|TYPE 2 DIAB WITH DIAB MCLR EDEMA, RESOLVED FOL TRTMT, UNSP
C2857155|T037|S72.111B|ICD10CM|DISPLACED FRACTURE OF GREATER TROCHANTER OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF GREATER TROCHANTER OF R FEMR, 7THB
C2857156|T037|S72.111C|ICD10CM|DISPLACED FRACTURE OF GREATER TROCHANTER OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF GREATER TROCHANTER OF R FEMR, 7THC
C2857154|T037|S72.111A|ICD10CM|DISPLACED FRACTURE OF GREATER TROCHANTER OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF GREATER TROCHANTER OF RIGHT FEMUR, INIT
C2857513|T037|S72.144A|ICD10CM|NONDISPLACED INTERTROCHANTERIC FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED INTERTROCHANTERIC FRACTURE OF RIGHT FEMUR, INIT
C2857514|T037|S72.144B|ICD10CM|NONDISPLACED INTERTROCHANTERIC FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP INTERTROCH FX RIGHT FEMUR, INIT FOR OPN FX TYPE I/2
C2857515|T037|S72.144C|ICD10CM|NONDISPLACED INTERTROCHANTERIC FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP INTERTROCH FX R FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2890022|T037|T82.518A|ICD10CM|BREAKDOWN (MECHANICAL) OF OTHER CARDIAC AND VASCULAR DEVICES AND IMPLANTS, INITIAL ENCOUNTER|BREAKDOWN OF CARDIAC AND VASCULAR DEVICES AND IMPLANTS, INIT
C2833941|T037|S14.126S|ICD10CM|CENTRAL CORD SYNDROME AT C6 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|CENTRAL CORD SYNDROME AT C6, SEQUELA
C2910920|T033|Z48.280|ICD10CM|ENCOUNTER FOR AFTERCARE FOLLOWING HEART-LUNG TRANSPLANT|ENCOUNTER FOR AFTERCARE FOLLOWING HEART-LUNG TRANSPLANT
C2833940|T037|S14.126D|ICD10CM|CENTRAL CORD SYNDROME AT C6 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|CENTRAL CORD SYNDROME AT C6, SUBS
C2901861|T047|M86.362|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, LEFT TIBIA AND FIBULA|CHRONIC MULTIFOCAL OSTEOMYELITIS, LEFT TIBIA AND FIBULA
C2833939|T037|S14.126A|ICD10CM|CENTRAL CORD SYNDROME AT C6 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|CENTRAL CORD SYNDROME AT C6, INIT
C2859231|T037|S73.036A|ICD10CM|OTHER ANTERIOR DISLOCATION OF UNSPECIFIED HIP, INITIAL ENCOUNTER|OTHER ANTERIOR DISLOCATION OF UNSPECIFIED HIP, INIT ENCNTR
C2901860|T047|M86.361|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, RIGHT TIBIA AND FIBULA|CHRONIC MULTIFOCAL OSTEOMYELITIS, RIGHT TIBIA AND FIBULA
C3251587|T046|T86.5|ICD10CM|COMPLICATIONS OF STEM CELL TRANSPLANT|COMPLICATIONS OF STEM CELL TRANSPLANT
C2901862|T047|M86.369|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, UNSPECIFIED TIBIA AND FIBULA|CHRONIC MULTIFOCAL OSTEOMYELITIS, UNSP TIBIA AND FIBULA
C2905689|T037|X73.8XXS|ICD10CM|INTENTIONAL SELF-HARM BY OTHER LARGER FIREARM DISCHARGE, SEQUELA|SELF-HARM BY OTH LARGER FIREARM DISCHARGE, SEQUELA
C2905687|T037|X73.8XXA|ICD10CM|INTENTIONAL SELF-HARM BY OTHER LARGER FIREARM DISCHARGE, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY OTH LARGER FIREARM DISCHARGE, INIT
C2856810|T037|S72.042A|ICD10CM|DISPLACED FRACTURE OF BASE OF NECK OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF BASE OF NECK OF LEFT FEMUR, INIT FOR CLOS FX
C2842133|T191|C50.829|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF UNSPECIFIED MALE BREAST|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF UNSP MALE BREAST
C2873940|T047|E08.638|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH OTHER ORAL COMPLICATIONS|DIABETES DUE TO UNDERLYING CONDITION W OTH ORAL COMP
C2856811|T037|S72.042B|ICD10CM|DISPLACED FRACTURE OF BASE OF NECK OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF BASE OF NECK OF L FEMUR, INIT FOR OPN FX TYPE I/2
C2842131|T191|C50.821|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF RIGHT MALE BREAST|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF RIGHT MALE BREAST
C2873939|T047|E08.630|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PERIODONTAL DISEASE|DIABETES DUE TO UNDERLYING CONDITION W PERIODONTAL DISEASE
C2832257|T037|S06.349A|ICD10CM|TRAUMATIC HEMORRHAGE OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|TRAUM HEMOR RIGHT CEREBRUM W LOC OF UNSP DURATION, INIT
C0236799|T048|F68.12|ICD10CM|FACTITIOUS DISORDER WITH PREDOMINANTLY PHYSICAL SIGNS AND SYMPTOMS|FACTITIOUS DISORDER W PREDOM PHYSICAL SIGNS AND SYMPTOMS
C0236798|T048|F68.13|ICD10CM|FACTITIOUS DISORDER WITH COMBINED PSYCHOLOGICAL AND PHYSICAL SIGNS AND SYMPTOMS|FACTITIOUS DISORD W COMB PSYCH AND PHYSCL SIGNS AND SYMPTOMS
C0015480|T048|F68.10|ICD10CM|FACTITIOUS DISORDER, UNSPECIFIED|FACTITIOUS DISORDER, UNSPECIFIED
C0015481|T048|F68.11|ICD10CM|FACTITIOUS DISORDER WITH PREDOMINANTLY PSYCHOLOGICAL SIGNS AND SYMPTOMS|FACTITIOUS DISORDER W PREDOM PSYCH SIGNS AND SYMPTOMS
C2832259|T037|S06.349S|ICD10CM|TRAUMATIC HEMORRHAGE OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|TRAUM HEMOR RIGHT CEREBRUM W LOC OF UNSP DURATION, SEQUELA
C2834058|T037|S14.157S|ICD10CM|OTHER INCOMPLETE LESION AT C7 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|OTH INCOMPLETE LESION AT C7, SEQUELA
C2883104|T047|I82.432|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF LEFT POPLITEAL VEIN|ACUTE EMBOLISM AND THROMBOSIS OF LEFT POPLITEAL VEIN
C2883105|T047|I82.433|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF POPLITEAL VEIN, BILATERAL|ACUTE EMBOLISM AND THROMBOSIS OF POPLITEAL VEIN, BILATERAL
C2873826|T047|D76.3|ICD10CM|OTHER HISTIOCYTOSIS SYNDROMES|RETICULOHISTIOCYTOMA (GIANT-CELL)
C2883103|T047|I82.431|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF RIGHT POPLITEAL VEIN|ACUTE EMBOLISM AND THROMBOSIS OF RIGHT POPLITEAL VEIN
C2874814|T048|F19.222|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE|OTH PSYCHOACTV SUBSTANCE DEPEND W INTOX W PERCEPTUAL DISTURB
C2874812|T048|F19.220|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH INTOXICATION, UNCOMPLICATED|OTH PSYCHOACTIVE SUBSTANCE DEPENDENCE W INTOXICATION, UNCOMP
C2883106|T047|I82.439|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED POPLITEAL VEIN|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED POPLITEAL VEIN
C2879799|T037|T47.5X2S|ICD10CM|POISONING BY DIGESTANTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY DIGESTANTS, INTENTIONAL SELF-HARM, SEQUELA
C2902730|T037|M96.629|ICD10CM|FRACTURE OF HUMERUS FOLLOWING INSERTION OF ORTHOPEDIC IMPLANT, JOINT PROSTHESIS, OR BONE PLATE, UNSPECIFIED ARM|FX HUMERUS FOL INSRT ORTHO IMPLNT/PROSTH/BONE PLT, UNSP ARM
C2889252|T047|M05.459|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSP HIP
C2890052|T037|T82.525A|ICD10CM|DISPLACEMENT OF UMBRELLA DEVICE, INITIAL ENCOUNTER|DISPLACEMENT OF UMBRELLA DEVICE, INITIAL ENCOUNTER
C2889250|T047|M05.451|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT HIP|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889251|T047|M05.452|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT HIP|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT HIP
C2889133|T047|M05.10|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP SITE
C4270598|T046|T85.735A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO CRANIAL OR SPINAL INFUSION CATHETER, INITIAL ENCOUNTER|I/I REACT D/T CRANIAL OR SPINAL INFUSION CATHETER, INIT
C3264025|T047|G43.829|ICD10CM|MENSTRUAL MIGRAINE, NOT INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|MENSTRUAL MIGRAINE, NOT INTRACTABLE, W/O STATUS MIGRAINOSUS
C2834057|T037|S14.157D|ICD10CM|OTHER INCOMPLETE LESION AT C7 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|OTH INCOMPLETE LESION AT C7, SUBS
C2869789|T037|S98.119A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED GREAT TOE, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF UNSP GREAT TOE, INIT ENCNTR
C2905660|T037|X71.3XXS|ICD10CM|INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION IN NATURAL WATER, SEQUELA|INTENTIONAL SELF-HARM BY DROWN IN NATURAL WATER, SEQUELA
C2858800|T037|S72.454B|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP SUPRCNDL FX W/O INTRCNDL EXTN LOW END R FEMR, 7THB
C2858801|T037|S72.454C|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP SUPRCNDL FX W/O INTRCNDL EXTN LOW END R FEMR, 7THC
C2902728|T037|M96.621|ICD10CM|FRACTURE OF HUMERUS FOLLOWING INSERTION OF ORTHOPEDIC IMPLANT, JOINT PROSTHESIS, OR BONE PLATE, RIGHT ARM|FX HUMERUS FOL INSRT ORTHO IMPLNT/PROSTH/BONE PLT, RIGHT ARM
C2890925|T037|T84.9XXA|ICD10CM|UNSPECIFIED COMPLICATION OF INTERNAL ORTHOPEDIC PROSTHETIC DEVICE, IMPLANT AND GRAFT, INITIAL ENCOUNTER|UNSP COMP OF INTERNAL ORTHOPEDIC PROSTH DEV/GRFT, INIT
C2858474|T037|S72.423A|ICD10CM|DISPLACED FRACTURE OF LATERAL CONDYLE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF LATERAL CONDYLE OF UNSP FEMUR, INIT FOR CLOS FX
C2838618|T037|S34.101S|ICD10CM|UNSPECIFIED INJURY TO L1 LEVEL OF LUMBAR SPINAL CORD, SEQUELA|UNSP INJURY TO L1 LEVEL OF LUMBAR SPINAL CORD, SEQUELA
C2858476|T037|S72.423C|ICD10CM|DISPLACED FRACTURE OF LATERAL CONDYLE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF LATERAL CONDYLE OF UNSP FEMR, 7THC
C2889324|T047|M05.679|ICD10CM|RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF UNSP ANK/FT W INVOLV OF ORGANS AND SYSTEMS
C2838617|T037|S34.101D|ICD10CM|UNSPECIFIED INJURY TO L1 LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY TO L1 LEVEL OF LUMBAR SPINAL CORD, SUBS ENCNTR
C2874387|T048|F10.229|ICD10CM|ALCOHOL DEPENDENCE WITH INTOXICATION, UNSPECIFIED|ALCOHOL DEPENDENCE WITH INTOXICATION, UNSPECIFIED
C2889322|T047|M05.671|ICD10CM|RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRIT OF RIGHT ANK/FT W INVOLV OF ORGANS AND SYSTEMS
C2889164|T047|M05.19|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS MULT SITE
C2874386|T048|F10.221|ICD10CM|ALCOHOL DEPENDENCE WITH INTOXICATION DELIRIUM|ALCOHOL DEPENDENCE WITH INTOXICATION DELIRIUM
C2874385|T048||ICD10CM|ALCOHOL DEPENDENCE WITH INTOXICATION, UNCOMPLICATED
C2842073|T191|C4A.72|ICD10CM|MERKEL CELL CARCINOMA OF LEFT LOWER LIMB, INCLUDING HIP|MERKEL CELL CARCINOMA OF LEFT LOWER LIMB, INCLUDING HIP
C2977926|T191|C4A.70|ICD10CM|MERKEL CELL CARCINOMA OF UNSPECIFIED LOWER LIMB, INCLUDING HIP|MERKEL CELL CARCINOMA OF UNSP LOWER LIMB, INCLUDING HIP
C2842072|T191|C4A.71|ICD10CM|MERKEL CELL CARCINOMA OF RIGHT LOWER LIMB, INCLUDING HIP|MERKEL CELL CARCINOMA OF RIGHT LOWER LIMB, INCLUDING HIP
C2876668|T037|T36.5X2A|ICD10CM|POISONING BY AMINOGLYCOSIDES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY AMINOGLYCOSIDES, INTENTIONAL SELF-HARM, INIT
C2859980|T037|S78.019D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT UNSPECIFIED HIP JOINT, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION AT UNSP HIP JOINT, SUBS ENCNTR
C2858320|T037|S72.409A|ICD10CM|UNSPECIFIED FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF LOWER END OF UNSP FEMUR, INIT FOR CLOS FX
C2858321|T037|S72.409B|ICD10CM|UNSPECIFIED FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP FX LOWER END OF UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2858322|T037|S72.409C|ICD10CM|UNSPECIFIED FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP FX LOWER END OF UNSP FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2876670|T037|T36.5X2S|ICD10CM|POISONING BY AMINOGLYCOSIDES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY AMINOGLYCOSIDES, INTENTIONAL SELF-HARM, SEQUELA
C2879870|T037|T47.8X2A|ICD10CM|POISONING BY OTHER AGENTS PRIMARILY AFFECTING GASTROINTESTINAL SYSTEM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH AGENTS AFF GI SYS, SELF-HARM, INIT
C2855865|T037|S68.110S|ICD10CM|COMPLETE TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF RIGHT INDEX FINGER, SEQUELA|COMPLETE TRAUMATIC MCP AMPUTATION OF R IDX FNGR, SEQUELA
C2838704|T037|S34.139D|ICD10CM|UNSPECIFIED INJURY TO SACRAL SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSPECIFIED INJURY TO SACRAL SPINAL CORD, SUBS ENCNTR
C2835254|T037|S22.029A|ICD10CM|UNSPECIFIED FRACTURE OF SECOND THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF SECOND THORACIC VERTEBRA, INIT FOR CLOS FX
C2835255|T037|S22.029B|ICD10CM|UNSPECIFIED FRACTURE OF SECOND THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF SECOND THORACIC VERTEBRA, INIT FOR OPN FX
C2857667|T037|S72.301A|ICD10CM|UNSPECIFIED FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF SHAFT OF RIGHT FEMUR, INIT FOR CLOS FX
C2857669|T037|S72.301C|ICD10CM|UNSPECIFIED FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP FX SHAFT OF RIGHT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2857668|T037|S72.301B|ICD10CM|UNSPECIFIED FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP FX SHAFT OF RIGHT FEMUR, INIT FOR OPN FX TYPE I/2
C2896566|T046|M80.049A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, UNSPECIFIED HAND, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, UNSP HAND, INIT
C2886208|T037|T65.92XA|ICD10CM|TOXIC EFFECT OF UNSPECIFIED SUBSTANCE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF UNSP SUBSTANCE, INTENTIONAL SELF-HARM, INIT
C2838703|T037|S34.139A|ICD10CM|UNSPECIFIED INJURY TO SACRAL SPINAL CORD, INITIAL ENCOUNTER|UNSPECIFIED INJURY TO SACRAL SPINAL CORD, INITIAL ENCOUNTER
C2874786|T048|F18.99|ICD10CM|INHALANT USE, UNSPECIFIED WITH UNSPECIFIED INHALANT-INDUCED DISORDER|INHALANT USE, UNSP WITH UNSP INHALANT-INDUCED DISORDER
C2889415|T047|M06.212|ICD10CM|RHEUMATOID BURSITIS, LEFT SHOULDER|RHEUMATOID BURSITIS, LEFT SHOULDER
C2884220|T037|T53.1X2S|ICD10CM|TOXIC EFFECT OF CHLOROFORM, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CHLOROFORM, INTENTIONAL SELF-HARM, SEQUELA
C2889414|T047|M06.211|ICD10CM|RHEUMATOID BURSITIS, RIGHT SHOULDER|RHEUMATOID BURSITIS, RIGHT SHOULDER
C2845927|T191|C69.92|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF LEFT EYE|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF LEFT EYE
C2845925|T191|C69.90|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF UNSPECIFIED EYE|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF UNSPECIFIED EYE
C2845926|T191|C69.91|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF RIGHT EYE|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF RIGHT EYE
C4237513|T048|F18.97|ICD10CM|INHALANT USE, UNSPECIFIED WITH INHALANT-INDUCED PERSISTING DEMENTIA|INHALANT-INDUCED MAJOR NEUROCOGNITIVE DISORDER
C4237567|T048|F18.94|ICD10CM|INHALANT USE, UNSPECIFIED WITH INHALANT-INDUCED MOOD DISORDER|INHALANT INDUCED DEPRESSIVE DISORDER
C4269405|T037|S02.40EA|ICD10CM|ZYGOMATIC FRACTURE, RIGHT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|ZYGOMATIC FRACTURE, RIGHT SIDE, INIT
C4269406|T037|S02.40EB|ICD10CM|ZYGOMATIC FRACTURE, RIGHT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|ZYGOMATIC FRACTURE, RIGHT SIDE, 7THB
C0342684|T047|E70.310|ICD10CM|X-LINKED OCULAR ALBINISM|X-LINKED OCULAR ALBINISM
C0268503|T019|E70.311|ICD10CM|AUTOSOMAL RECESSIVE OCULAR ALBINISM|AUTOSOMAL RECESSIVE OCULAR ALBINISM
C2874229|T019|E70.318|ICD10CM|OTHER OCULAR ALBINISM|OTHER OCULAR ALBINISM
C2874379|T048|F10.181|ICD10CM|ALCOHOL ABUSE WITH ALCOHOL-INDUCED SEXUAL DYSFUNCTION|ALCOHOL ABUSE WITH ALCOHOL-INDUCED SEXUAL DYSFUNCTION
C2838301|T037|S32.476B|ICD10CM|NONDISPLACED FRACTURE OF MEDIAL WALL OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP FX OF MEDIAL WALL OF UNSP ACETAB, INIT FOR OPN FX
C0838561|T047|M46.99|ICD10AM|UNSPECIFIED INFLAMMATORY SPONDYLOPATHY, MULTIPLE SITES IN SPINE|UNSPECIFIED INFLAMMATORY SPONDYLOPATHY, SITE UNSPECIFIED
C2833338|T037|S12.231A|ICD10CM|UNSPECIFIED TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP TRAUM NONDISP SPONDYLOLYSIS OF THIRD CERVCAL VERT, INIT
C4270403|T046|T83.722A|ICD10CM|EXPOSURE OF IMPLANTED URETHRAL MESH INTO URETHRA, INITIAL ENCOUNTER|EXPOSURE OF IMPLANTED URETHRAL MESH INTO URETHRA, INIT
C2876545|T037|T36.0X2A|ICD10CM|POISONING BY PENICILLINS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY PENICILLINS, INTENTIONAL SELF-HARM, INIT ENCNTR
C2889464|T046|M06.379|ICD10CM|RHEUMATOID NODULE, UNSPECIFIED ANKLE AND FOOT|RHEUMATOID NODULE, UNSPECIFIED ANKLE AND FOOT
C0838560|T047|M46.98|ICD10CM|UNSPECIFIED INFLAMMATORY SPONDYLOPATHY, SACRAL AND SACROCOCCYGEAL REGION|UNSP INFLAMMATORY SPONDYLOPATHY, SACR/SACROCYGL REGION
C2889462|T046|M06.371|ICD10CM|RHEUMATOID NODULE, RIGHT ANKLE AND FOOT|RHEUMATOID NODULE, RIGHT ANKLE AND FOOT
C2889463|T046|M06.372|ICD10CM|RHEUMATOID NODULE, LEFT ANKLE AND FOOT|RHEUMATOID NODULE, LEFT ANKLE AND FOOT
C0349023|T191|C47.4|DMDICD10|MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF ABDOMEN|BOESARTIGE NEUBILDUNG: PERIPHERE NERVEN DES ABDOMENS
C0349024|T191|C47.5|DMDICD10|MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF PELVIS|BOESARTIGE NEUBILDUNG: PERIPHERE NERVEN DES BECKENS
C2977921|T191|C47.6|ICD10CM|MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF TRUNK, UNSPECIFIED|MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF UNSPECIFIED PART OF TRUNK
C0349019|T191|C47.0|DMDICD10|MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF HEAD, FACE AND NECK|BOESARTIGE NEUBILDUNG: PERIPHERE NERVEN DES KOPFES, DES GESICHTES UND DES HALSES
C0349022|T191|C47.3|DMDICD10|MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF THORAX|BOESARTIGE NEUBILDUNG: PERIPHERE NERVEN DES THORAX
C0348358|T191|C47.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF PERIPHERAL NERVES AND AUTONOMIC NERVOUS SYSTEM|BOESARTIGE NEUBILDUNG: PERIPHERE NERVEN UND AUTONOMES NERVENSYSTEM, MEHRERE TEILBEREICHE UEBERLAPPEND
C2977922|T191|C47.9|ICD10CM|MALIGNANT NEOPLASM OF PERIPHERAL NERVES AND AUTONOMIC NERVOUS SYSTEM, UNSPECIFIED|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF PERIPHERAL NERVES AND AUTONOMIC NERVOUS SYSTEM
C2890784|T037|T84.420A|ICD10CM|DISPLACEMENT OF MUSCLE AND TENDON GRAFT, INITIAL ENCOUNTER|DISPLACEMENT OF MUSCLE AND TENDON GRAFT, INITIAL ENCOUNTER
C2857428|T037|S72.135A|ICD10CM|NONDISPLACED APOPHYSEAL FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED APOPHYSEAL FRACTURE OF LEFT FEMUR, INIT
C2832323|T037|S06.364S|ICD10CM|TRAUMATIC HEMORRHAGE OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|TRAUM HEMOR CEREB, W LOC OF 6 HOURS TO 24 HOURS, SEQUELA
C2874979|T048|F63.89|ICD10CM|OTHER IMPULSE DISORDERS|OTHER IMPULSE DISORDERS
C2832321|T037|S06.364A|ICD10CM|TRAUMATIC HEMORRHAGE OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|TRAUM HEMOR CEREB, W LOC OF 6 HOURS TO 24 HOURS, INIT
C0021776|T048||ICD10CM|INTERMITTENT EXPLOSIVE DISORDER
C2890563|T037|T84.092A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTERNAL RIGHT KNEE PROSTHESIS, INITIAL ENCOUNTER|MECH COMPL OF INTERNAL RIGHT KNEE PROSTHESIS, INIT ENCNTR
C2876207|T037|T32.65|ICD10CM|CORROSIONS INVOLVING 60-69% OF BODY SURFACE WITH 50-59% THIRD DEGREE CORROSION|CORROS 60-69% OF BODY SURFACE W 50-59% THIRD DEGREE CORROS
C0010481|T047|E24.9|DMDICD10|CUSHING'S SYNDROME, UNSPECIFIED|CUSHING-SYNDROM, NICHT NAEHER BEZEICHNET
C0348458|T047|E24.8|DMDICD10|OTHER CUSHING'S SYNDROME|SONSTIGES CUSHING-SYNDROM
C2890634|T037|T84.124A|ICD10CM|DISPLACEMENT OF INTERNAL FIXATION DEVICE OF RIGHT FEMUR, INITIAL ENCOUNTER|DISPLACEMENT OF INT FIX OF RIGHT FEMUR, INIT
C0342446|T047|E24.4|DMDICD10|ALCOHOL-INDUCED PSEUDO-CUSHING'S SYNDROME|ALKOHOLINDUZIERTES PSEUDO-CUSHING-SYNDROM
C0027577|T191|E24.1|DMDICD10|NELSON'S SYNDROME|NELSON-TUMOR
C0342712|T047|E71.2|DMDICD10|DISORDER OF BRANCHED-CHAIN AMINO-ACID METABOLISM, UNSPECIFIED|STOERUNG DES STOFFWECHSELS VERZWEIGTER AMINOSAEUREN, NICHT NAEHER BEZEICHNET
C0001231|T047|E24.3|DMDICD10|ECTOPIC ACTH SYNDROME|EKTOPISCHES ACTH-SYNDROM
C3714740|T047|E24.2|DMDICD10|DRUG-INDUCED CUSHING'S SYNDROME|ARZNEIMITTELINDUZIERTES CUSHING-SYNDROM
C2889995|T037|T82.49XD|ICD10CM|OTHER COMPLICATION OF VASCULAR DIALYSIS CATHETER, SUBSEQUENT ENCOUNTER|OTH COMPLICATION OF VASCULAR DIALYSIS CATHETER, SUBS ENCNTR
C2869902|T037|S98.921S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT FOOT, LEVEL UNSPECIFIED, SEQUELA|PARTIAL TRAUMATIC AMP OF RIGHT FOOT, LEVEL UNSP, SEQUELA
C2901906|T047|M86.559|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED FEMUR|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED FEMUR
C2837926|T037|S32.413A|ICD10CM|DISPLACED FRACTURE OF ANTERIOR WALL OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF ANTERIOR WALL OF UNSP ACETABULUM, INIT
C2832348|T037|S06.370S|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF CEREBELLUM WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|CONTUS/LAC/HEM CRBLM W/O LOSS OF CONSCIOUSNESS, SEQUELA
C2901904|T047|M86.551|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, RIGHT FEMUR|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, RIGHT FEMUR
C2877867|T037|T41.0X2A|ICD10CM|POISONING BY INHALED ANESTHETICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY INHALED ANESTHETICS, SELF-HARM, INIT
C2901905|T047|M86.552|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, LEFT FEMUR|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, LEFT FEMUR
C2869900|T037|S98.921A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT FOOT, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF RIGHT FOOT, LEVEL UNSP, INIT
C2832346|T037|S06.370A|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF CEREBELLUM WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|CONTUS/LAC/HEM CRBLM W/O LOSS OF CONSCIOUSNESS, INIT
C2877869|T037|T41.0X2S|ICD10CM|POISONING BY INHALED ANESTHETICS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY INHALED ANESTHETICS, SELF-HARM, SEQUELA
C2848408|T037|S58.022S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT ELBOW LEVEL, LEFT ARM, SEQUELA|PARTIAL TRAUMATIC AMP AT ELBOW LEVEL, LEFT ARM, SEQUELA
C4270581|T046|T85.732A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO IMPLANTED ELECTRONIC NEUROSTIMULATOR OF PERIPHERAL NERVE, ELECTRODE (LEAD), INITIAL ENCOUNTER|I/I REACT D/T IMPLNT ELEC NSTIM OF PRPH NRV, LEAD, INIT
C2882085|T047|I13.11|ICD10CM|HYPERTENSIVE HEART AND CHRONIC KIDNEY DISEASE WITHOUT HEART FAILURE, WITH STAGE 5 CHRONIC KIDNEY DISEASE, OR END STAGE RENAL DISEASE|HYP HRT AND CHR KDNY DIS W/O HRT FAIL, W STG 5 CHR KDNY/ESRD
C2882084|T047|I13.10|ICD10CM|HYPERTENSIVE HEART AND CHRONIC KIDNEY DISEASE WITHOUT HEART FAILURE, WITH STAGE 1 THROUGH STAGE 4 CHRONIC KIDNEY DISEASE, OR UNSPECIFIED CHRONIC KIDNEY DISEASE|HYP HRT & CHR KDNY DIS W/O HRT FAIL, W STG 1-4/UNSP CHR KDNY
C0854199|T191||ICD10CM|CHRONIC MYELOMONOCYTIC LEUKEMIA, IN REMISSION
C2861620|T191|C93.10|ICD10CM|CHRONIC MYELOMONOCYTIC LEUKEMIA NOT HAVING ACHIEVED REMISSION|CHRONIC MYELOMONOCYTIC LEUKEMIA NOT ACHIEVE REMISSION
C2848406|T037|S58.022A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT ELBOW LEVEL, LEFT ARM, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION AT ELBOW LEVEL, LEFT ARM, INIT
C2366868|T191||ICD10CM|CHRONIC MYELOMONOCYTIC LEUKEMIA, IN RELAPSE
C2882397|T047|I63.49|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF OTHER CEREBRAL ARTERY|CEREBRAL INFARCTION DUE TO EMBOLISM OF OTHER CEREBRAL ARTERY
C2833993|T037|S14.141A|ICD10CM|BROWN-SEQUARD SYNDROME AT C1 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|BROWN-SEQUARD SYNDROME AT C1, INIT
C2833189|T037|S12.041A|ICD10CM|NONDISPLACED LATERAL MASS FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP LATERAL MASS FX FIRST CERVCAL VERTEBRA, INIT
C2857017|T037|S72.065B|ICD10CM|NONDISPLACED ARTICULAR FRACTURE OF HEAD OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP ARTIC FX HEAD OF L FEMUR, INIT FOR OPN FX TYPE I/2
C2857018|T037|S72.065C|ICD10CM|NONDISPLACED ARTICULAR FRACTURE OF HEAD OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP ARTIC FX HEAD OF L FEMR, INIT FOR OPN FX TYPE 3A/B/C
C2855949|T037|S68.411S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT HAND AT WRIST LEVEL, SEQUELA|COMPLETE TRAUMATIC AMP OF RIGHT HAND AT WRIST LEVEL, SEQUELA
C2882380|T047|I63.40|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF UNSPECIFIED CEREBRAL ARTERY|CEREBRAL INFARCTION DUE TO EMBOLISM OF UNSP CEREBRAL ARTERY
C3264378|T047|I67.841|ICD10CM|REVERSIBLE CEREBROVASCULAR VASOCONSTRICTION SYNDROME|REVERSIBLE CEREBROVASCULAR VASOCONSTRICTION SYNDROME
C3264379|T047|I67.848|ICD10CM|OTHER CEREBROVASCULAR VASOSPASM AND VASOCONSTRICTION|OTHER CEREBROVASCULAR VASOSPASM AND VASOCONSTRICTION
C2833986|T037|S14.138S|ICD10CM|ANTERIOR CORD SYNDROME AT C8 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|ANTERIOR CORD SYNDROME AT C8, SEQUELA
C2877441|T037|T39.312S|ICD10CM|POISONING BY PROPIONIC ACID DERIVATIVES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY PROPIONIC ACID DERIVATIVES, SELF-HARM, SEQUELA
C2885835|T037|T63.712S|ICD10CM|TOXIC EFFECT OF CONTACT WITH VENOMOUS MARINE PLANT, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CNTCT W VENOM MARINE PLANT, SLF-HRM, SEQUELA
C2833984|T037|S14.138A|ICD10CM|ANTERIOR CORD SYNDROME AT C8 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|ANTERIOR CORD SYNDROME AT C8, INIT
C2877439|T037|T39.312A|ICD10CM|POISONING BY PROPIONIC ACID DERIVATIVES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY PROPIONIC ACID DERIVATIVES, SELF-HARM, INIT
C2885833|T037|T63.712A|ICD10CM|TOXIC EFFECT OF CONTACT WITH VENOMOUS MARINE PLANT, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CONTACT W VENOM MARINE PLANT, SLF-HRM, INIT
C2833985|T037|S14.138D|ICD10CM|ANTERIOR CORD SYNDROME AT C8 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|ANTERIOR CORD SYNDROME AT C8, SUBS
C2876190|T037|T32.33|ICD10CM|CORROSIONS INVOLVING 30-39% OF BODY SURFACE WITH 30-39% THIRD DEGREE CORROSION|CORROS 30-39% OF BODY SURFACE W 30-39% THIRD DEGREE CORROS
C2876189|T037|T32.32|ICD10CM|CORROSIONS INVOLVING 30-39% OF BODY SURFACE WITH 20-29% THIRD DEGREE CORROSION|CORROS 30-39% OF BODY SURFACE W 20-29% THIRD DEGREE CORROS
C2876188|T037|T32.31|ICD10CM|CORROSIONS INVOLVING 30-39% OF BODY SURFACE WITH 10-19% THIRD DEGREE CORROSION|CORROS 30-39% OF BODY SURFACE W 10-19% THIRD DEGREE CORROS
C2501076|T060|B410|ICD10PCS|PULMONARY PARACOCCIDIOIDOMYCOSIS|IMAGING @ LOWER ARTERIES @ FLUOROSCOPY @ ABDOMINAL AORTA
C2889379|T047|M05.869|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED KNEE|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSP KNEE
C2889377|T047|M05.861|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT KNEE|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF RIGHT KNEE
C2889378|T047|M05.862|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT KNEE|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT KNEE
C2833870|T037|S14.107A|ICD10CM|UNSPECIFIED INJURY AT C7 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY AT C7 LEVEL OF CERVICAL SPINAL CORD, INIT ENCNTR
C2833871|T037|S14.107D|ICD10CM|UNSPECIFIED INJURY AT C7 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY AT C7 LEVEL OF CERVICAL SPINAL CORD, SUBS ENCNTR
C2833872|T037|S14.107S|ICD10CM|UNSPECIFIED INJURY AT C7 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|UNSP INJURY AT C7 LEVEL OF CERVICAL SPINAL CORD, SEQUELA
C1279420|T048||ICD10CM|GENERALIZED ANXIETY DISORDER
C0086769|T048||ICD10CM|PANIC DISORDER [EPISODIC PAROXYSMAL ANXIETY]
C2838670|T037|S34.122A|ICD10CM|INCOMPLETE LESION OF L2 LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|INCOMPLETE LESION OF L2 LEVEL OF LUMBAR SPINAL CORD, INIT
C2838671|T037|S34.122D|ICD10CM|INCOMPLETE LESION OF L2 LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|INCOMPLETE LESION OF L2 LEVEL OF LUMBAR SPINAL CORD, SUBS
C0838554|T047|M46.92|ICD10AM|UNSPECIFIED INFLAMMATORY SPONDYLOPATHY, CERVICAL REGION|UNSPECIFIED INFLAMMATORY SPONDYLOPATHY, CERVICAL REGION
C2893629|T047|M12.011|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], RIGHT SHOULDER|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], RIGHT SHOULDER
C0041657|T033||ICD10CM|UNSPECIFIED COMA
C2832523|T037|S06.6X3S|ICD10CM|TRAUMATIC SUBARACHNOID HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, SEQUELA|TRAUM SUBRAC HEM W LOC OF 1-5 HRS 59 MIN, SEQUELA
C2977074|T047|J96.91|ICD10CM|RESPIRATORY FAILURE, UNSPECIFIED WITH HYPOXIA|RESPIRATORY FAILURE, UNSPECIFIED WITH HYPOXIA
C2977073|T047|J96.90|ICD10CM|RESPIRATORY FAILURE, UNSPECIFIED, UNSPECIFIED WHETHER WITH HYPOXIA OR HYPERCAPNIA|RESPIRATORY FAILURE, UNSP, UNSP W HYPOXIA OR HYPERCAPNIA
C2977075|T047|J96.92|ICD10CM|RESPIRATORY FAILURE, UNSPECIFIED WITH HYPERCAPNIA|RESPIRATORY FAILURE, UNSPECIFIED WITH HYPERCAPNIA
C2860142|T037|S79.111A|ICD10CM|SALTER-HARRIS TYPE I PHYSEAL FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SLTR-HARIS TYPE I PHYSEAL FX LOWER END OF RIGHT FEMUR, INIT
C2832521|T037|S06.6X3A|ICD10CM|TRAUMATIC SUBARACHNOID HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|TRAUM SUBRAC HEM W LOC OF 1-5 HRS 59 MIN, INIT
C2885491|T037|T63.192A|ICD10CM|TOXIC EFFECT OF VENOM OF OTHER REPTILES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF REPTILES, SELF-HARM, INIT
C2882753|T047|I70.312|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, LEFT LEG|ATHSCL UNSP TYPE BYPASS OF EXTRM W INTRMT CLAUD, LEFT LEG
C2889180|T047|M05.241|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT HAND|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889181|T047|M05.242|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT HAND|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT HAND
C2882752|T047|I70.311|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, RIGHT LEG|ATHSCL UNSP TYPE BYPASS OF EXTRM W INTRMT CLAUD, RIGHT LEG
C2889179|T047|M05.249|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND
C2882755|T047|I70.318|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, OTHER EXTREMITY|ATHSCL UNSP TYPE BYPASS OF EXTRM W INTRMT CLAUD, OTH EXTRM
C2882756|T047|I70.319|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, UNSPECIFIED EXTREMITY|ATHSCL UNSP TYPE BYPASS OF EXTRM W INTRMT CLAUD, UNSP EXTRM
C2874592|T048|F14.221|ICD10CM|COCAINE DEPENDENCE WITH INTOXICATION DELIRIUM|COCAINE DEPENDENCE WITH INTOXICATION DELIRIUM
C2874591|T048||ICD10CM|COCAINE DEPENDENCE WITH INTOXICATION, UNCOMPLICATED
C2874593|T048|F14.222|ICD10CM|COCAINE DEPENDENCE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE|COCAINE DEPENDENCE W INTOXICATION W PERCEPTUAL DISTURBANCE
C2835773|T037|S24.109D|ICD10CM|UNSPECIFIED INJURY AT UNSPECIFIED LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY AT UNSP LEVEL OF THORACIC SPINAL CORD, SUBS
C2887830|T047|K51.80|ICD10CM|OTHER ULCERATIVE COLITIS WITHOUT COMPLICATIONS|OTHER ULCERATIVE COLITIS WITHOUT COMPLICATIONS
C2883310|T037|T49.1X2S|ICD10CM|POISONING BY ANTIPRURITICS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ANTIPRURITICS, INTENTIONAL SELF-HARM, SEQUELA
C2837803|T037|S32.301A|ICD10CM|UNSPECIFIED FRACTURE OF RIGHT ILIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF RIGHT ILIUM, INIT FOR CLOS FX
C2837804|T037|S32.301B|ICD10CM|UNSPECIFIED FRACTURE OF RIGHT ILIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF RIGHT ILIUM, INIT ENCNTR FOR OPEN FRACTURE
C2832635|T037|S06.891A|ICD10CM|OTHER SPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|INTCRAN INJ W LOC OF 30 MINUTES OR LESS, INIT
C4237397|T048|F13.921|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH INTOXICATION DELIRIUM|SEDATIVE, HYPNOTIC, OR ANXIOLYTIC-INDUCED DELIRIUM
C2874553|T048|F13.920|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH INTOXICATION, UNCOMPLICATED|SEDATV/HYP/ANXIOLYTC USE, UNSP W INTOXICATION, UNCOMPLICATED
C2874541|T048|F13.251|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|SEDATV/HYP/ANXIOLYTC DEPEND W PSYCHOTIC DISORDER W HALLUCIN
C2874540|T048|F13.250|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|SEDATV/HYP/ANXIOLYTC DEPEND W PSYCHOTIC DISORDER W DELUSIONS
C2858697|T037|S72.444C|ICD10CM|NONDISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF LOW EPIPHY (SEPARATION) OF R FEMR, 7THC
C2874555|T048|F13.929|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH INTOXICATION, UNSPECIFIED|SEDATV/HYP/ANXIOLYTC USE, UNSP W INTOXICATION, UNSP
C2874542|T048|F13.25|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED PSYCHOTIC DISORDER
C2900881|T046|M84.419A|ICD10CM|PATHOLOGICAL FRACTURE, UNSPECIFIED SHOULDER, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, UNSP SHOULDER, INIT FOR FX
C2879621|T037|T46.902S|ICD10CM|POISONING BY UNSPECIFIED AGENTS PRIMARILY AFFECTING THE CARDIOVASCULAR SYSTEM, INTENTIONAL SELF-HARM, SEQUELA|POISN BY UNSP AGENTS AFF THE CARDIOVASC SYS, SLF-HRM, SQLA
C4268781|T046|M84.755A|ICD10CM|COMPLETE TRANSVERSE ATYPICAL FEMORAL FRACTURE, LEFT LEG, INITIAL ENCOUNTER FOR FRACTURE|COMPLETE TRANSVERSE ATYP FEMORAL FRACTURE, LEFT LEG, INIT
C2835176|T037|S22.008B|ICD10CM|OTHER FRACTURE OF UNSPECIFIED THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF UNSP THORACIC VERTEBRA, INIT FOR OPN FX
C2879619|T037|T46.902A|ICD10CM|POISONING BY UNSPECIFIED AGENTS PRIMARILY AFFECTING THE CARDIOVASCULAR SYSTEM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY UNSP AGENTS AFF THE CARDIOVASC SYS, SELF-HARM, INIT
C0153474|T191|C31.9|DMDICD10|MALIGNANT NEOPLASM OF ACCESSORY SINUS, UNSPECIFIED|BOESARTIGE NEUBILDUNG: NASENNEBENHOEHLE, NICHT NAEHER BEZEICHNET
C0349041|T191|C31.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF ACCESSORY SINUSES|BOESARTIGE NEUBILDUNG: NASENNEBENHOEHLEN, MEHRERE TEILBEREICHE UEBERLAPPEND
C2882841|T047|I70.449|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF UNSPECIFIED SITE|ATHSCL AUTOL VEIN BYPASS OF LEFT LEG W ULCER OF UNSP SITE
C2845891|T191|C64.9|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED KIDNEY, EXCEPT RENAL PELVIS|MALIGNANT NEOPLASM OF UNSP KIDNEY, EXCEPT RENAL PELVIS
C0153477|T191|C31.1|DMDICD10|MALIGNANT NEOPLASM OF ETHMOIDAL SINUS|BOESARTIGE NEUBILDUNG: SINUS ETHMOIDALIS [SIEBBEINZELLEN]
C2837943|T191|C31.0|ICD10CM|MALIGNANT NEOPLASM OF MAXILLARY SINUS|MALIGNANT NEOPLASM OF ANTRUM (HIGHMORE) (MAXILLARY)
C0153479|T191|C31.3|DMDICD10|MALIGNANT NEOPLASM OF SPHENOID SINUS|BOESARTIGE NEUBILDUNG: SINUS SPHENOIDALIS [KEILBEINHOEHLE]
C0153478|T191|C31.2|DMDICD10|MALIGNANT NEOPLASM OF FRONTAL SINUS|BOESARTIGE NEUBILDUNG: SINUS FRONTALIS [STIRNHOEHLE]
C2977941|T191|C64.2|ICD10CM|MALIGNANT NEOPLASM OF LEFT KIDNEY, EXCEPT RENAL PELVIS|MALIGNANT NEOPLASM OF LEFT KIDNEY, EXCEPT RENAL PELVIS
C2845890|T191|C64.1|ICD10CM|MALIGNANT NEOPLASM OF RIGHT KIDNEY, EXCEPT RENAL PELVIS|MALIGNANT NEOPLASM OF RIGHT KIDNEY, EXCEPT RENAL PELVIS
C3263998|T047|G40.B01|ICD10CM|JUVENILE MYOCLONIC EPILEPSY, NOT INTRACTABLE, WITH STATUS EPILEPTICUS|JUVENILE MYOCLONIC EPILEPSY, NOT INTRACTABLE, W STAT EPI
C2901942|T046|M87.029|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED HUMERUS|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED HUMERUS
C2879568|T037|T46.7X2A|ICD10CM|POISONING BY PERIPHERAL VASODILATORS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY PERIPHERAL VASODILATORS, SELF-HARM, INIT
C3263999|T047|G40.B09|ICD10CM|JUVENILE MYOCLONIC EPILEPSY, NOT INTRACTABLE, WITHOUT STATUS EPILEPTICUS|JUVENILE MYOCLONIC EPILEPSY, NOT INTRACTABLE, W/O STAT EPI
C2901940|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF RIGHT HUMERUS
C2902362|T047|M89.619|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, UNSPECIFIED SHOULDER|OSTEOPATHY AFTER POLIOMYELITIS, UNSPECIFIED SHOULDER
C2876176|T037|T31.94|ICD10CM|BURNS INVOLVING 90% OR MORE OF BODY SURFACE WITH 40-49% THIRD DEGREE BURNS|BURNS OF 90%/MORE OF BODY SURFC W 40-49% THIRD DEGREE BURNS
C2902361|T047|M89.612|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, LEFT SHOULDER|OSTEOPATHY AFTER POLIOMYELITIS, LEFT SHOULDER
C2902360|T047|M89.611|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, RIGHT SHOULDER|OSTEOPATHY AFTER POLIOMYELITIS, RIGHT SHOULDER
C2876177|T037|T31.95|ICD10CM|BURNS INVOLVING 90% OR MORE OF BODY SURFACE WITH 50-59% THIRD DEGREE BURNS|BURNS OF 90%/MORE OF BODY SURFC W 50-59% THIRD DEGREE BURNS
C2712603|T056||ICD9CM|IODINE-DEFICIENCY RELATED DIFFUSE (ENDEMIC) GOITER
C2873858|T047|E01.1|ICD10CM|IODINE-DEFICIENCY RELATED MULTINODULAR (ENDEMIC) GOITER|IODINE-DEFICIENCY RELATED NODULAR GOITER
C2712624|T056|E012|ICD9CM|IODINE-DEFICIENCY RELATED (ENDEMIC) GOITER, UNSPECIFIED|ACTIVITIES INVOLVING ARTS AND HANDCRAFTS
C4269286|T037|S02.11BA|ICD10CM|TYPE I OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE I OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, INIT
C2712943|T056|E018|ICD9CM|OTHER IODINE-DEFICIENCY RELATED THYROID DISORDERS AND ALLIED CONDITIONS|ACTIVITIES INVOLVING PLAYING MUSICAL INSTRUMENT
C2876180|T037|T31.98|ICD10CM|BURNS INVOLVING 90% OR MORE OF BODY SURFACE WITH 80-89% THIRD DEGREE BURNS|BURNS OF 90%/MORE OF BODY SURFC W 80-89% THIRD DEGREE BURNS
C2876181|T037|T31.99|ICD10CM|BURNS INVOLVING 90% OR MORE OF BODY SURFACE WITH 90% OR MORE THIRD DEGREE BURNS|BURNS OF 90%/MORE OF BODY SURFC W 90%/MORE THIRD DEG BURNS
C2910940|T033|Z49.02|ICD10CM|ENCOUNTER FOR FITTING AND ADJUSTMENT OF PERITONEAL DIALYSIS CATHETER|ENCOUNTER FOR FIT/ADJST OF PERITONEAL DIALYSIS CATHETER
C2910939|T033|Z49.01|ICD10CM|ENCOUNTER FOR FITTING AND ADJUSTMENT OF EXTRACORPOREAL DIALYSIS CATHETER|ENCOUNTER FOR FITTING AND ADJUSTMENT OF EXTRACORPOREAL DIALYSIS CATHETER
C2883482|T037|T49.8X2A|ICD10CM|POISONING BY OTHER TOPICAL AGENTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH TOPICAL AGENTS, INTENTIONAL SELF-HARM, INIT
C2857737|T037|S72.322B|ICD10CM|DISPLACED TRANSVERSE FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL TRANSVERSE FX SHAFT OF L FEMR, 7THB
C2857738|T037|S72.322C|ICD10CM|DISPLACED TRANSVERSE FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL TRANSVERSE FX SHAFT OF L FEMR, 7THC
C2857736|T037|S72.322A|ICD10CM|DISPLACED TRANSVERSE FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED TRANSVERSE FRACTURE OF SHAFT OF LEFT FEMUR, INIT
C2875351|T047|G83.24|ICD10CM|MONOPLEGIA OF UPPER LIMB AFFECTING LEFT NONDOMINANT SIDE|MONOPLEGIA OF UPPER LIMB AFFECTING LEFT NONDOMINANT SIDE
C2875350|T047|G83.23|ICD10CM|MONOPLEGIA OF UPPER LIMB AFFECTING RIGHT NONDOMINANT SIDE|MONOPLEGIA OF UPPER LIMB AFFECTING RIGHT NONDOMINANT SIDE
C2875349|T047|G83.22|ICD10CM|MONOPLEGIA OF UPPER LIMB AFFECTING LEFT DOMINANT SIDE|MONOPLEGIA OF UPPER LIMB AFFECTING LEFT DOMINANT SIDE
C2875348|T047|G83.21|ICD10CM|MONOPLEGIA OF UPPER LIMB AFFECTING RIGHT DOMINANT SIDE|MONOPLEGIA OF UPPER LIMB AFFECTING RIGHT DOMINANT SIDE
C0154703|T047|G83.2|ICD10CM|MONOPLEGIA OF UPPER LIMB AFFECTING UNSPECIFIED SIDE|MONOPLEGIA OF UPPER LIMB
C2857035|T037|S72.066C|ICD10CM|NONDISPLACED ARTICULAR FRACTURE OF HEAD OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP ARTIC FX HEAD OF UNSP FEMR, 7THC
C2875378|T047|G90.59|ICD10CM|COMPLEX REGIONAL PAIN SYNDROME I OF OTHER SPECIFIED SITE|COMPLEX REGIONAL PAIN SYNDROME I OF OTHER SPECIFIED SITE
C2859972|T037|S78.011D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT RIGHT HIP JOINT, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION AT RIGHT HIP JOINT, SUBS
C2857033|T037|S72.066A|ICD10CM|NONDISPLACED ARTICULAR FRACTURE OF HEAD OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED ARTICULAR FRACTURE OF HEAD OF UNSP FEMUR, INIT
C2875367|T047|G90.5|ICD10CM|COMPLEX REGIONAL PAIN SYNDROME I, UNSPECIFIED|COMPLEX REGIONAL PAIN SYNDROME I (CRPS I)
C0339946|T047|A21.2|DMDICD10|PULMONARY TULAREMIA|PULMONALE TULARAEMIE
C2838122|T037|S32.435B|ICD10CM|NONDISPLACED FRACTURE OF ANTERIOR COLUMN [ILIOPUBIC] OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP FX OF ANT COLUMN OF LEFT ACETAB, INIT FOR OPN FX
C2838121|T037|S32.435A|ICD10CM|NONDISPLACED FRACTURE OF ANTERIOR COLUMN [ILIOPUBIC] OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF ANTERIOR COLUMN OF LEFT ACETABULUM, INIT
C2859973|T037|S78.011S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT RIGHT HIP JOINT, SEQUELA|COMPLETE TRAUMATIC AMPUTATION AT RIGHT HIP JOINT, SEQUELA
C2837488|T037|S32.011A|ICD10CM|STABLE BURST FRACTURE OF FIRST LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|STABLE BURST FRACTURE OF FIRST LUMBAR VERTEBRA, INIT
C2837489|T037|S32.011B|ICD10CM|STABLE BURST FRACTURE OF FIRST LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|STABLE BURST FRACTURE OF FIRST LUM VERTEBRA, INIT FOR OPN FX
C2878537|T037|T43.592S|ICD10CM|POISONING BY OTHER ANTIPSYCHOTICS AND NEUROLEPTICS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH ANTIPSYCHOT/NEUROLEPT, SELF-HARM, SEQUELA
C1579029|T047||ICD10CM|CHRONIC KIDNEY DISEASE, UNSPECIFIED
C2316810|T047|N18.6|ICD10CM|END STAGE RENAL DISEASE|END STAGE RENAL DISEASE
C2316810|T047|N18.6|ICD10CM|CHRONIC KIDNEY DISEASE, STAGE 5|END STAGE RENAL DISEASE
C1561641|T047|N18.4|ICD10CM|CHRONIC KIDNEY DISEASE, STAGE 4 (SEVERE)|CHRONIC KIDNEY DISEASE, STAGE 4 (SEVERE)
C1561640|T047|N18.3|ICD10CM|CHRONIC KIDNEY DISEASE, STAGE 3 (MODERATE)|CHRONIC KIDNEY DISEASE, STAGE 3 (MODERATE)
C1561639|T047|N18.2|ICD10CM|CHRONIC KIDNEY DISEASE, STAGE 2 (MILD)|CHRONIC KIDNEY DISEASE, STAGE 2 (MILD)
C2316401|T047||ICD10CM|CHRONIC KIDNEY DISEASE, STAGE 1
C2856053|T037|S68.622S|ICD10CM|PARTIAL TRAUMATIC TRANSPHALANGEAL AMPUTATION OF RIGHT MIDDLE FINGER, SEQUELA|PARTIAL TRAUMATIC TRNSPHAL AMP OF R MID FINGER, SEQUELA
C2878535|T037|T43.592A|ICD10CM|POISONING BY OTHER ANTIPSYCHOTICS AND NEUROLEPTICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH ANTIPSYCHOT/NEUROLEPT, SELF-HARM, INIT
C0522624|T191|C86.3|ICD10CM|SUBCUTANEOUS PANNICULITIS-LIKE T-CELL LYMPHOMA|SUBCUTANEOUS PANNICULITIS-LIKE T-CELL LYMPHOMA
C2854066|T191|C86.2|ICD10CM|ENTEROPATHY-TYPE (INTESTINAL) T-CELL LYMPHOMA|ENTEROPATHY-TYPE (INTESTINAL) T-CELL LYMPHOMA
C2854065|T047|C86.1|ICD10CM|HEPATOSPLENIC T-CELL LYMPHOMA|ALPHA-BETA AND GAMMA DELTA TYPES
C0392788|T191||ICD10CM|EXTRANODAL NK/T-CELL LYMPHOMA, NASAL TYPE
C2854068|T191|C86.6|ICD10CM|PRIMARY CUTANEOUS CD30-POSITIVE T-CELL PROLIFERATIONS|PRIMARY CUTANEOUS CD30-POSITIVE T-CELL PROLIFERATIONS
C0020981|T191|C86.5|ICD10CM|ANGIOIMMUNOBLASTIC T-CELL LYMPHOMA|ANGIOIMMUNOBLASTIC T-CELL LYMPHOMA
C4509017|T191|C86.4|ICD10CM|BLASTIC NK-CELL LYMPHOMA|BLASTIC PLASMACYTOID DENDRITIC CELL NEOPLASM (BPDCN)
C0339966|T047|J18.1|ICD10CM|LOBAR PNEUMONIA, UNSPECIFIED ORGANISM|LOBAR PNEUMONIA, UNSPECIFIED ORGANISM
C2889898|T037|T82.311A|ICD10CM|BREAKDOWN (MECHANICAL) OF CAROTID ARTERIAL GRAFT (BYPASS), INITIAL ENCOUNTER|BREAKDOWN OF CAROTID ARTERIAL GRAFT (BYPASS), INIT
C2901328|T046|M84.573A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, UNSPECIFIED ANKLE, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, UNSP ANKLE, INIT
C2877489|T037|T39.4X2S|ICD10CM|POISONING BY ANTIRHEUMATICS, NOT ELSEWHERE CLASSIFIED, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ANTIRHEUMATICS, NEC, SELF-HARM, SEQUELA
C2857548|T037|S72.146B|ICD10CM|NONDISPLACED INTERTROCHANTERIC FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP INTERTROCH FX UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2857549|T037|S72.146C|ICD10CM|NONDISPLACED INTERTROCHANTERIC FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP INTERTROCH FX UNSP FEMR, INIT FOR OPN FX TYPE 3A/B/C
C2857547|T037|S72.146A|ICD10CM|NONDISPLACED INTERTROCHANTERIC FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED INTERTROCHANTERIC FRACTURE OF UNSP FEMUR, INIT
C2885091|T037|T60.8X2A|ICD10CM|TOXIC EFFECT OF OTHER PESTICIDES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF OTH PESTICIDES, INTENTIONAL SELF-HARM, INIT
C2877487|T037|T39.4X2A|ICD10CM|POISONING BY ANTIRHEUMATICS, NOT ELSEWHERE CLASSIFIED, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ANTIRHEUMATICS, NEC, SELF-HARM, INIT
C2885093|T037|T60.8X2S|ICD10CM|TOXIC EFFECT OF OTHER PESTICIDES, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF PESTICIDES, INTENTIONAL SELF-HARM, SEQUELA
C0838494|T047|M46.02|ICD10AM|SPINAL ENTHESOPATHY, CERVICAL REGION|SPINAL ENTHESOPATHY, CERVICAL REGION
C0838495|T047|M46.03|ICD10AM|SPINAL ENTHESOPATHY, CERVICOTHORACIC REGION|SPINAL ENTHESOPATHY, CERVICOTHORACIC REGION
C0838492|T047|M46.00|ICD10AM|SPINAL ENTHESOPATHY, SITE UNSPECIFIED|SPINAL ENTHESOPATHY, MULTIPLE SITES IN SPINE
C0838493|T047|M46.01|ICD10AM|SPINAL ENTHESOPATHY, OCCIPITO-ATLANTO-AXIAL REGION|SPINAL ENTHESOPATHY, OCCIPITO-ATLANTO-AXIAL REGION
C0838498|T047|M46.06|ICD10AM|SPINAL ENTHESOPATHY, LUMBAR REGION|SPINAL ENTHESOPATHY, LUMBAR REGION
C0838499|T047|M46.07|ICD10AM|SPINAL ENTHESOPATHY, LUMBOSACRAL REGION|SPINAL ENTHESOPATHY, LUMBOSACRAL REGION
C0838496|T047|M46.04|ICD10AM|SPINAL ENTHESOPATHY, THORACIC REGION|SPINAL ENTHESOPATHY, THORACIC REGION
C0838497|T047|M46.05|ICD10AM|SPINAL ENTHESOPATHY, THORACOLUMBAR REGION|SPINAL ENTHESOPATHY, THORACOLUMBAR REGION
C0838500|T047|M46.08|ICD10AM|SPINAL ENTHESOPATHY, SACRAL AND SACROCOCCYGEAL REGION|SPINAL ENTHESOPATHY, SACRAL AND SACROCOCCYGEAL REGION
C0838492|T047|M46.09|ICD10CM|SPINAL ENTHESOPATHY, MULTIPLE SITES IN SPINE|SPINAL ENTHESOPATHY, MULTIPLE SITES IN SPINE
C2854038|T191|C85.25|ICD10CM|MEDIASTINAL (THYMIC) LARGE B-CELL LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|MEDIASTNL LG B-CELL LYMPH, NODES OF ING RGN AND LOWER LIMB
C2853844|T191|C82.56|ICD10CM|DIFFUSE FOLLICLE CENTER LYMPHOMA, INTRAPELVIC LYMPH NODES|DIFFUSE FOLLICLE CENTER LYMPHOMA, INTRAPELVIC LYMPH NODES
C2854040|T191|C85.27|ICD10CM|MEDIASTINAL (THYMIC) LARGE B-CELL LYMPHOMA, SPLEEN|MEDIASTINAL (THYMIC) LARGE B-CELL LYMPHOMA, SPLEEN
C2854039|T191|C85.26|ICD10CM|MEDIASTINAL (THYMIC) LARGE B-CELL LYMPHOMA, INTRAPELVIC LYMPH NODES|MEDIASTINAL (THYMIC) LARGE B-CELL LYMPHOMA, INTRAPELV NODES
C2854034|T191|C85.21|ICD10CM|MEDIASTINAL (THYMIC) LARGE B-CELL LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK|MEDIASTNL LARGE B-CELL LYMPH, NODES OF HEAD, FACE, AND NECK
C0742803|T047||ICD10CM|CONUS MEDULLARIS SYNDROME
C2854036|T191|C85.23|ICD10CM|MEDIASTINAL (THYMIC) LARGE B-CELL LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES|MEDIASTINAL (THYMIC) LARGE B-CELL LYMPHOMA, INTRA-ABD NODES
C2854035|T191|C85.22|ICD10CM|MEDIASTINAL (THYMIC) LARGE B-CELL LYMPHOMA, INTRATHORACIC LYMPH NODES|MEDIASTNL (THYMIC) LARGE B-CELL LYMPHOMA, INTRATHORAC NODES
C4270495|T046|T85.190A|ICD10CM|OTHER MECHANICAL COMPLICATION OF IMPLANTED ELECTRONIC NEUROSTIMULATOR OF BRAIN ELECTRODE (LEAD), INITIAL ENCOUNTER|MECH COMPL OF IMPLNT ELEC NSTIM OF BRAIN LEAD, INIT
C2854042|T191|C85.29|ICD10CM|MEDIASTINAL (THYMIC) LARGE B-CELL LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES|MEDIASTNL LARGE B-CELL LYMPH, EXTRNOD AND SOLID ORGAN SITES
C0477423|T047|G95.8|ICD10CM|OTHER SPECIFIED DISEASES OF SPINAL CORD|OTHER SPECIFIED DISEASES OF SPINAL CORD
C2853847|T191|C82.59|ICD10CM|DIFFUSE FOLLICLE CENTER LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES|DIFFUSE FOLICL CENTER LYMPH, EXTRNOD AND SOLID ORGAN SITES
C2853846|T191|C82.58|ICD10CM|DIFFUSE FOLLICLE CENTER LYMPHOMA, LYMPH NODES OF MULTIPLE SITES|DIFFUSE FOLLICLE CENTER LYMPHOMA, LYMPH NODES MULT SITE
C0342261|T047|E10.69|ICD10AM|TYPE 1 DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATION|TYPE 1 DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATION
C2902039|T046|M87.222|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, LEFT HUMERUS|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, LEFT HUMERUS
C2874070|T047||ICD10CM|TYPE 1 DIABETES MELLITUS WITH HYPERGLYCEMIA
C2876203|T037|T32.61|ICD10CM|CORROSIONS INVOLVING 60-69% OF BODY SURFACE WITH 10-19% THIRD DEGREE CORROSION|CORROS 60-69% OF BODY SURFACE W 10-19% THIRD DEGREE CORROS
C1535090|T047|I27.81|ICD10CM|COR PULMONALE (CHRONIC)|COR PULMONALE (CHRONIC)
C4509221|T047|I27.83|ICD10CM|EISENMENGER'S SYNDROME|PULMONARY HYPERTENSION WITH RIGHT TO LEFT SHUNT RELATED TO CONGENITAL HEART DISEASE
C0856722|T046|I27.82|ICD10CM|CHRONIC PULMONARY EMBOLISM|CHRONIC PULMONARY EMBOLISM
C0348595|T047|I27.89|ICD10CM|OTHER SPECIFIED PULMONARY HEART DISEASES|OTHER SPECIFIED PULMONARY HEART DISEASES
C2832385|T037|S06.379S|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF CEREBELLUM WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|CONTUS/LAC/HEM CRBLM W LOC OF UNSP DURATION, SEQUELA
C2902040|T046|M87.229|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED HUMERUS|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED HUMERUS
C1328840|T047|D89.82|ICD10CM|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME [ALPS]|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME [ALPS]
C2860120|T037|S79.101A|ICD10CM|UNSPECIFIED PHYSEAL FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP PHYSEAL FRACTURE OF LOWER END OF RIGHT FEMUR, INIT
C0869046|T047|D89.89|ICD10CM|OTHER SPECIFIED DISORDERS INVOLVING THE IMMUNE MECHANISM, NOT ELSEWHERE CLASSIFIED|OTH DISRD INVOLVING THE IMMUNE MECHANISM, NEC
C2876204|T037|T32.62|ICD10CM|CORROSIONS INVOLVING 60-69% OF BODY SURFACE WITH 20-29% THIRD DEGREE CORROSION|CORROS 60-69% OF BODY SURFACE W 20-29% THIRD DEGREE CORROS
C2856673|T037|S72.026C|ICD10CM|NONDISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF EPIPHY (SEPARATION) (UPPER) OF UNSP FEMR, 7THC
C2900555|T046|M80.872A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, LEFT ANKLE AND FOOT, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, LEFT ANK/FT, INIT
C2859223|T037|S73.034A|ICD10CM|OTHER ANTERIOR DISLOCATION OF RIGHT HIP, INITIAL ENCOUNTER|OTHER ANTERIOR DISLOCATION OF RIGHT HIP, INITIAL ENCOUNTER
C2901852|T047|M86.341|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, RIGHT HAND|CHRONIC MULTIFOCAL OSTEOMYELITIS, RIGHT HAND
C2901853|T047|M86.342|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, LEFT HAND|CHRONIC MULTIFOCAL OSTEOMYELITIS, LEFT HAND
C2901854|T047|M86.349|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, UNSPECIFIED HAND|CHRONIC MULTIFOCAL OSTEOMYELITIS, UNSPECIFIED HAND
C2833932|T037|S14.124D|ICD10CM|CENTRAL CORD SYNDROME AT C4 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|CENTRAL CORD SYNDROME AT C4, SUBS
C2833931|T037|S14.124A|ICD10CM|CENTRAL CORD SYNDROME AT C4 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|CENTRAL CORD SYNDROME AT C4, INIT
C2873757|T033|D56.2|ICD10CM|DELTA-BETA THALASSEMIA|HOMOZYGOUS DELTA-BETA THALASSEMIA
C2873756|T047||ICD10CM|BETA THALASSEMIA
C3161175|T047|D56.0|ICD10CM|ALPHA THALASSEMIA|HYDROPS FETALIS DUE TO ALPHA THALASSEMIA
C2882632|T047|I69.859|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING UNSPECIFIED SIDE|HEMIPLGA FOLLOWING OTH CEREBVASC DISEASE AFFECTING UNSP SIDE
C0019025|T047|D56.4|DMDICD10|HEREDITARY PERSISTENCE OF FETAL HEMOGLOBIN [HPFH]|HEREDITAERE PERSISTENZ FETALEN HAEMOGLOBINS [HPFH]
C2831484|T037|S02.411A|ICD10CM|LEFORT I FRACTURE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|LEFORT I FRACTURE, INITIAL ENCOUNTER FOR CLOSED FRACTURE
C2831485|T037|S02.411B|ICD10CM|LEFORT I FRACTURE, INITIAL ENCOUNTER FOR OPEN FRACTURE|LEFORT I FRACTURE, INITIAL ENCOUNTER FOR OPEN FRACTURE
C2882631|T047|I69.854|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING LEFT NON-DOMINANT SIDE|HEMIPLGA FOL OTH CEREBVASC DISEASE AFF LEFT NONDOM SIDE
C2882630|T047|I69.853|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING RIGHT NON-DOMINANT SIDE|HEMIPLGA FOL OTH CEREBVASC DISEASE AFF RIGHT NONDOM SIDE
C2882629|T047|I69.852|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING LEFT DOMINANT SIDE|HEMIPLGA FOL OTH CEREBVASC DISEASE AFF LEFT DOMINANT SIDE
C2882628|T047|I69.851|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING RIGHT DOMINANT SIDE|HEMIPLGA FOL OTH CEREBVASC DISEASE AFF RIGHT DOMINANT SIDE
C2873931|T047|E08.618|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH OTHER DIABETIC ARTHROPATHY|DIABETES DUE TO UNDERLYING CONDITION W OTH DIABETIC ARTHROP
C2842114|T191|C50.519|ICD10CM|MALIGNANT NEOPLASM OF LOWER-OUTER QUADRANT OF UNSPECIFIED FEMALE BREAST|MALIG NEOPLASM OF LOWER-OUTER QUADRANT OF UNSP FEMALE BREAST
C2873930|T047|E08.610|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH DIABETIC NEUROPATHIC ARTHROPATHY|DIABETES DUE TO UNDRL COND W DIABETIC NEUROPATHIC ARTHROP
C2842112|T191|C50.511|ICD10CM|MALIGNANT NEOPLASM OF LOWER-OUTER QUADRANT OF RIGHT FEMALE BREAST|MALIG NEOPLM OF LOWER-OUTER QUADRANT OF RIGHT FEMALE BREAST
C2842113|T191|C50.512|ICD10CM|MALIGNANT NEOPLASM OF LOWER-OUTER QUADRANT OF LEFT FEMALE BREAST|MALIG NEOPLASM OF LOWER-OUTER QUADRANT OF LEFT FEMALE BREAST
C2831489|T037|S02.411S|ICD10CM|LEFORT I FRACTURE, SEQUELA|LEFORT I FRACTURE, SEQUELA
C2833360|T037|S12.251A|ICD10CM|OTHER TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH TRAUM NONDISP SPONDYLOLYSIS OF THIRD CERVCAL VERT, INIT
C2890036|T037|T82.521A|ICD10CM|DISPLACEMENT OF SURGICALLY CREATED ARTERIOVENOUS SHUNT, INITIAL ENCOUNTER|DISPLACEMENT OF SURGICALLY CREATED ARTERIOVENOUS SHUNT, INIT
C2833361|T037|S12.251B|ICD10CM|OTHER TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH TRAUM NONDISP SPONDYLOLYSIS OF 3RD CERVCAL VERT, 7THB
C2857085|T037|S72.099A|ICD10CM|OTHER FRACTURE OF HEAD AND NECK OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF HEAD AND NECK OF UNSP FEMUR, INIT
C4509316|T047|L97.518|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF RIGHT FOOT WITH OTHER SPECIFIED SEVERITY|NON-PRS CHRONIC ULCER OTH PRT RIGHT FOOT WITH OTH SEVERITY
C2888727|T047|L97.519|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF RIGHT FOOT WITH UNSPECIFIED SEVERITY|NON-PRS CHRONIC ULCER OTH PRT RIGHT FOOT W UNSP SEVERITY
C2888726|T047|L97.514|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF RIGHT FOOT WITH NECROSIS OF BONE|NON-PRS CHRONIC ULCER OTH PRT RIGHT FOOT W NECROSIS OF BONE
C4509314|T047|L97.515|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF RIGHT FOOT WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OTH PRT R FOOT WITH MSL INVL W/O EVD OF NECR
C4509315|T047|L97.516|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF RIGHT FOOT WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OTH PRT R FOOT WITH BNE INVL W/O EVD OF NECR
C2888723|T047|L97.511|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF RIGHT FOOT LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHRONIC ULCER OTH PRT R FOOT LIMITED TO BRKDWN SKIN
C2888724|T047|L97.512|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF RIGHT FOOT WITH FAT LAYER EXPOSED|NON-PRS CHRONIC ULCER OTH PRT RIGHT FOOT W FAT LAYER EXPOSED
C2888725|T047|L97.513|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF RIGHT FOOT WITH NECROSIS OF MUSCLE|NON-PRS CHRONIC ULCER OTH PRT RIGHT FOOT W NECROS MUSCLE
C2874671|T048|F15.950|ICD10CM|OTHER STIMULANT USE, UNSPECIFIED WITH STIMULANT-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|OTH STIM USE, UNSP W STIM-INDUCE PSYCH DISORDER W DELUSIONS
C2874672|T048|F15.951|ICD10CM|OTHER STIMULANT USE, UNSPECIFIED WITH STIMULANT-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|OTH STIM USE, UNSP W STIM-INDUCE PSYCH DISORDER W HALLUCIN
C2889260|T047|M05.472|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF LEFT ANK/FT
C2889259|T047|M05.471|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF RIGHT ANK/FT
C4236974|T048|F15.959|ICD10CM|OTHER STIMULANT USE, UNSPECIFIED WITH STIMULANT-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|AMPHETAMINE OR OTHER STIMULANT-INDUCED PSYCHOTIC DISORDER, WITHOUT USE DISORDER
C2883093|T047|I82.411|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF RIGHT FEMORAL VEIN|ACUTE EMBOLISM AND THROMBOSIS OF RIGHT FEMORAL VEIN
C2889261|T047|M05.479|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF UNSP ANK/FT
C2883095|T047|I82.413|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF FEMORAL VEIN, BILATERAL|ACUTE EMBOLISM AND THROMBOSIS OF FEMORAL VEIN, BILATERAL
C2856605|T037|S72.022C|ICD10CM|DISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF EPIPHY (SEPARATION) (UPPER) OF L FEMR, 7THC
C2856604|T037|S72.022B|ICD10CM|DISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF EPIPHY (SEPARATION) (UPPER) OF L FEMR, 7THB
C2856603|T037|S72.022A|ICD10CM|DISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF EPIPHYSIS (SEPARATION) (UPPER) OF L FEMUR, INIT
C2835342|T037|S22.051B|ICD10CM|STABLE BURST FRACTURE OF T5-T6 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|STABLE BURST FRACTURE OF T5-T6 VERTEBRA, INIT FOR OPN FX
C1135210|T047|I77.79|ICD10CM|DISSECTION OF OTHER SPECIFIED ARTERY|DISSECTION OF OTHER SPECIFIED ARTERY
C2835341|T037|S22.051A|ICD10CM|STABLE BURST FRACTURE OF T5-T6 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|STABLE BURST FRACTURE OF T5-T6 VERTEBRA, INIT FOR CLOS FX
C4268550|T047||ICD10CM|DISSECTION OF ARTERY OF LOWER EXTREMITY
C4076498|T047|I77.76|ICD10CM|DISSECTION OF ARTERY OF UPPER EXTREMITY|DISSECTION OF ARTERY OF UPPER EXTREMITY
C4270822|T047|I77.75|ICD10CM|DISSECTION OF OTHER PRECEREBRAL ARTERIES|DISSECTION OF BASILAR ARTERY (TRUNK)
C0338586|T047||ICD10CM|DISSECTION OF VERTEBRAL ARTERY
C0919563|T047|I77.73|ICD10CM|DISSECTION OF RENAL ARTERY|DISSECTION OF RENAL ARTERY
C0340649|T047|I77.72|ICD10CM|DISSECTION OF ILIAC ARTERY|DISSECTION OF ILIAC ARTERY
C0338585|T047|I77.71|ICD10CM|DISSECTION OF CAROTID ARTERY|DISSECTION OF CAROTID ARTERY
C4268548|T047|I77.70|ICD10CM|DISSECTION OF UNSPECIFIED ARTERY|DISSECTION OF UNSPECIFIED ARTERY
C2878252|T037|T42.8X2A|ICD10CM|POISONING BY ANTIPARKINSONISM DRUGS AND OTHER CENTRAL MUSCLE-TONE DEPRESSANTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY ANTIPARKNS DRUG/CENTR MUSC-TONE DEPR, SLF-HRM, INIT
C0001916|T047|E70.30|ICD10CM|ALBINISM, UNSPECIFIED|ALBINISM, UNSPECIFIED
C2857087|T037|S72.099C|ICD10CM|OTHER FRACTURE OF HEAD AND NECK OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|OTH FX HEAD/NECK OF UNSP FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2874233|T019|E70.39|ICD10CM|OTHER SPECIFIED ALBINISM|OTHER SPECIFIED ALBINISM
C4268085|T047|E11.3412|ICD10CM|TYPE 2 DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|TYPE 2 DIAB WITH SEVERE NONP RTNOP WITH MACULAR EDEMA, L EYE
C4268086|T047|E11.3413|ICD10CM|TYPE 2 DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|TYPE 2 DIAB WITH SEVERE NONP RTNOP WITH MACULAR EDEMA, BI
C2874274|T047|E75.29|ICD10CM|OTHER SPHINGOLIPIDOSIS|FARBER'S SYNDROME
C2901249|T046|M84.551A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, RIGHT FEMUR, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, RIGHT FEMUR, INIT
C2890854|T037|T84.619A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL FIXATION DEVICE OF UNSPECIFIED BONE OF ARM, INITIAL ENCOUNTER|INFECT/INFLM REACT DUE TO INT FIX OF UNSP BONE OF ARM, INIT
C2833331|T037|S12.230A|ICD10CM|UNSPECIFIED TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP TRAUM DISPL SPONDYLOLYSIS OF THIRD CERVCAL VERT, INIT
C0017205|T047||ICD10CM|GAUCHER DISEASE
C0023521|T047||ICD10CM|KRABBE DISEASE
C2833384|T037|S12.300B|ICD10CM|UNSPECIFIED DISPLACED FRACTURE OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP DISP FX OF FOURTH CERVICAL VERTEBRA, INIT FOR OPN FX
C0002986|T047||ICD10CM|FABRY (-ANDERSON) DISEASE
C4269567|T037|S02.80XB|ICD10CM|FRACTURE OF OTHER SPECIFIED SKULL AND FACIAL BONES, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FX OTH SKULL AND FACIAL BONES, UNSPECIFIED SIDE, 7THB
C2833332|T037|S12.230B|ICD10CM|UNSPECIFIED TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP TRAUM DISPL SPONDYLOLYSIS OF 3RD CERVCAL VERT, 7THB
C0023522|T047||ICD10CM|METACHROMATIC LEUKODYSTROPHY
C2845874|T191|C62.02|ICD10CM|MALIGNANT NEOPLASM OF UNDESCENDED LEFT TESTIS|MALIGNANT NEOPLASM OF UNDESCENDED LEFT TESTIS
C2889315|T047|M05.652|ICD10CM|RHEUMATOID ARTHRITIS OF LEFT HIP WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF LEFT HIP W INVOLV OF ORGANS AND SYSTEMS
C2889314|T047|M05.651|ICD10CM|RHEUMATOID ARTHRITIS OF RIGHT HIP WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF RIGHT HIP W INVOLV OF ORGANS AND SYSTEMS
C2845873|T191|C62.01|ICD10CM|MALIGNANT NEOPLASM OF UNDESCENDED RIGHT TESTIS|MALIGNANT NEOPLASM OF UNDESCENDED RIGHT TESTIS
C2882909|T047|I70.591|ICD10CM|OTHER ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, RIGHT LEG|OTH ATHSCL NONAUT BIO BYPASS OF THE EXTREMITIES, RIGHT LEG
C2889316|T047|M05.659|ICD10CM|RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF UNSP HIP W INVOLV OF ORGANS AND SYSTEMS
C2900860|T046|M84.40XA|ICD10CM|PATHOLOGICAL FRACTURE, UNSPECIFIED SITE, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, UNSP SITE, INIT ENCNTR FOR FRACTURE
C2858441|T037|S72.421B|ICD10CM|DISPLACED FRACTURE OF LATERAL CONDYLE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF LATERAL CONDYLE OF R FEMR, 7THB
C2858442|T037|S72.421C|ICD10CM|DISPLACED FRACTURE OF LATERAL CONDYLE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF LATERAL CONDYLE OF R FEMR, 7THC
C2835240|T037|S22.022A|ICD10CM|UNSTABLE BURST FRACTURE OF SECOND THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSTABLE BURST FRACTURE OF SECOND THORACIC VERTEBRA, INIT
C2835241|T037|S22.022B|ICD10CM|UNSTABLE BURST FRACTURE OF SECOND THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSTABLE BURST FX SECOND THOR VERTEBRA, INIT FOR OPN FX
C2877464|T037|T39.392S|ICD10CM|POISONING BY OTHER NONSTEROIDAL ANTI-INFLAMMATORY DRUGS [NSAID], INTENTIONAL SELF-HARM, SEQUELA|POISN BY OTH NONSTEROID ANTI-INFLAM DRUGS, SLF-HRM, SEQUELA
C2843334|T037|S48.921A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT SHOULDER AND UPPER ARM, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|PARTIAL TRAUM AMP OF RIGHT SHLDR/UP ARM, LEVEL UNSP, INIT
C2886750|T037|T79.A0XA|ICD10CM|COMPARTMENT SYNDROME, UNSPECIFIED, INITIAL ENCOUNTER|COMPARTMENT SYNDROME, UNSPECIFIED, INITIAL ENCOUNTER
C2843336|T037|S48.921S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT SHOULDER AND UPPER ARM, LEVEL UNSPECIFIED, SEQUELA|PARTIAL TRAUM AMP OF RIGHT SHLDR/UP ARM, LEVEL UNSP, SEQUELA
C2882913|T047|I70.599|ICD10CM|OTHER ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, UNSPECIFIED EXTREMITY|OTH ATHSCL NONAUT BIO BYPASS OF THE EXTRM, UNSP EXTREMITY
C2874299|T047|E83.19|ICD10CM|OTHER DISORDERS OF IRON METABOLISM|OTHER DISORDERS OF IRON METABOLISM
C2884498|T037|T56.2X2S|ICD10CM|TOXIC EFFECT OF CHROMIUM AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CHROMIUM AND ITS COMPND, SELF-HARM, SEQUELA
C2883073|T047|I80.232|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF LEFT TIBIAL VEIN|PHLEBITIS AND THROMBOPHLEBITIS OF LEFT TIBIAL VEIN
C2883074|T047|I80.233|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF TIBIAL VEIN, BILATERAL|PHLEBITIS AND THROMBOPHLEBITIS OF TIBIAL VEIN, BILATERAL
C2977008|T047|I82.5Y1|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF RIGHT PROXIMAL LOWER EXTREMITY|CHR EMBLSM AND THOMBOS UNSP DEEP VEINS OF R PROX LOW EXTRM
C2884496|T037|T56.2X2A|ICD10CM|TOXIC EFFECT OF CHROMIUM AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CHROMIUM AND ITS COMPOUNDS, SELF-HARM, INIT
C0348829|T047|J95.1|DMDICD10|ACUTE PULMONARY INSUFFICIENCY FOLLOWING THORACIC SURGERY|AKUTE PULMONALE INSUFFIZIENZ NACH THORAXOPERATION
C0348830|T047|J95.2|DMDICD10|ACUTE PULMONARY INSUFFICIENCY FOLLOWING NONTHORACIC SURGERY|AKUTE PULMONALE INSUFFIZIENZ NACH NICHT AM THORAX VORGENOMMENER OPERATION
C0348831|T047|J95.3|DMDICD10|CHRONIC PULMONARY INSUFFICIENCY FOLLOWING SURGERY|CHRONISCHE PULMONALE INSUFFIZIENZ NACH OPERATION
C2855873|T037|S68.112S|ICD10CM|COMPLETE TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF RIGHT MIDDLE FINGER, SEQUELA|COMPLETE TRAUMATIC MCP AMPUTATION OF R MID FINGER, SEQUELA
C2884482|T037|T56.1X2S|ICD10CM|TOXIC EFFECT OF MERCURY AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF MERCURY AND ITS COMPND, SELF-HARM, SEQUELA
C2902062|T046|M87.256|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED FEMUR|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED FEMUR
C2902060|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, RIGHT FEMUR
C2902059|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, PELVIS
C2902061|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, LEFT FEMUR
C0839938|T047|M86.19|ICD10CM|OTHER ACUTE OSTEOMYELITIS, MULTIPLE SITES|OTHER ACUTE OSTEOMYELITIS, MULTIPLE SITES
C2837960|T191|C34.90|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED PART OF UNSPECIFIED BRONCHUS OR LUNG|MALIGNANT NEOPLASM OF UNSP PART OF UNSP BRONCHUS OR LUNG
C2837961|T191|C34.91|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED PART OF RIGHT BRONCHUS OR LUNG|MALIGNANT NEOPLASM OF UNSP PART OF RIGHT BRONCHUS OR LUNG
C2837962|T191|C34.92|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED PART OF LEFT BRONCHUS OR LUNG|MALIGNANT NEOPLASM OF UNSP PART OF LEFT BRONCHUS OR LUNG
C0348587|T047|I15.1|DMDICD10|HYPERTENSION SECONDARY TO OTHER RENAL DISORDERS|HYPERTONIE ALS FOLGE VON SONSTIGEN NIERENKRANKHEITEN
C0020545|T047|I15.0|DMDICD10|RENOVASCULAR HYPERTENSION|RENOVASKULAERE HYPERTONIE
C2882781|T047|I70.344|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF HEEL AND MIDFOOT|ATHSCL UNSP TYPE BYPASS OF LEFT LEG W ULC OF HEEL AND MIDFT
C0155616|T047|I15|DMDICD10|SECONDARY HYPERTENSION, UNSPECIFIED|SEKUNDAERE HYPERTONIE
C0348586|T047|I15.8|DMDICD10|OTHER SECONDARY HYPERTENSION|SONSTIGE SEKUNDAERE HYPERTONIE
C2889421|T047|M06.231|ICD10CM|RHEUMATOID BURSITIS, RIGHT WRIST|RHEUMATOID BURSITIS, RIGHT WRIST
C2889422|T047|M06.232|ICD10CM|RHEUMATOID BURSITIS, LEFT WRIST|RHEUMATOID BURSITIS, LEFT WRIST
C4269396|T037|S02.40CS|ICD10CM|MAXILLARY FRACTURE, RIGHT SIDE, SEQUELA|MAXILLARY FRACTURE, RIGHT SIDE, SEQUELA
C2889423|T047|M06.239|ICD10CM|RHEUMATOID BURSITIS, UNSPECIFIED WRIST|RHEUMATOID BURSITIS, UNSPECIFIED WRIST
C0007965|T047|D72.0|ICD10CM|CHEDIAK-HIGASHI SYNDROME|HEREDITARY LEUKOMELANOPATHY
C0079504|T047||ICD10CM|HERMANSKY-PUDLAK SYNDROME
C2842064|T191|C4A.52|ICD10CM|MERKEL CELL CARCINOMA OF SKIN OF BREAST|MERKEL CELL CARCINOMA OF SKIN OF BREAST
C0152486|T047|A02.1|DMDICD10|SALMONELLA SEPSIS|SALMONELLENSEPSIS
C2874232|T019|E70.338|ICD10CM|OTHER ALBINISM WITH HEMATOLOGIC ABNORMALITY|OTHER ALBINISM WITH HEMATOLOGIC ABNORMALITY
C2874231|T019|E70.339|ICD10CM|ALBINISM WITH HEMATOLOGIC ABNORMALITY, UNSPECIFIED|ALBINISM WITH HEMATOLOGIC ABNORMALITY, UNSPECIFIED
C4269391|T037|S02.40CA|ICD10CM|MAXILLARY FRACTURE, RIGHT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|MAXILLARY FRACTURE, RIGHT SIDE, INIT
C2877843|T037|T40.992S|ICD10CM|POISONING BY OTHER PSYCHODYSLEPTICS [HALLUCINOGENS], INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH PSYCHODYSLEPTICS, SELF-HARM, SEQUELA
C2879644|T037|T46.992A|ICD10CM|POISONING BY OTHER AGENTS PRIMARILY AFFECTING THE CARDIOVASCULAR SYSTEM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY OTH AGENTS AFF THE CARDIOVASC SYS, SELF-HARM, INIT
C2890441|T037|T84.023A|ICD10CM|INSTABILITY OF INTERNAL LEFT KNEE PROSTHESIS, INITIAL ENCOUNTER|INSTABILITY OF INTERNAL LEFT KNEE PROSTHESIS, INIT ENCNTR
C2877841|T037|T40.992A|ICD10CM|POISONING BY OTHER PSYCHODYSLEPTICS [HALLUCINOGENS], INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH PSYCHODYSLEPTICS, SELF-HARM, INIT
C2889456|T046|M06.352|ICD10CM|RHEUMATOID NODULE, LEFT HIP|RHEUMATOID NODULE, LEFT HIP
C2889455|T046|M06.351|ICD10CM|RHEUMATOID NODULE, RIGHT HIP|RHEUMATOID NODULE, RIGHT HIP
C2896706|T046|M80.831A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, RIGHT FOREARM, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, R FOREARM, INIT
C0264511|T047|J84.2|ICD10CM|LYMPHOID INTERSTITIAL PNEUMONIA|LYMPHOID INTERSTITIAL PNEUMONIA
C2889457|T046|M06.359|ICD10CM|RHEUMATOID NODULE, UNSPECIFIED HIP|RHEUMATOID NODULE, UNSPECIFIED HIP
C2900997|T046|M84.452A|ICD10CM|PATHOLOGICAL FRACTURE, LEFT FEMUR, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, LEFT FEMUR, INIT ENCNTR FOR FRACTURE
C2843310|T037|S48.121S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN RIGHT SHOULDER AND ELBOW, SEQUELA|PARTIAL TRAUM AMP AT LEVEL BETW R SHLDR AND ELBOW, SEQUELA
C2885223|T037|T62.0X2S|ICD10CM|TOXIC EFFECT OF INGESTED MUSHROOMS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF INGESTED MUSHROOMS, SELF-HARM, SEQUELA
C0346110|T191|C45.2|DMDICD10|MESOTHELIOMA OF PERICARDIUM|MESOTHELIOM DES PERIKARDS
C0812413|T191|C45.0|DMDICD10|MESOTHELIOMA OF PLEURA|MESOTHELIOM DER PLEURA
C3714724|T191|C45.1|ICD10CM|MESOTHELIOMA OF PERITONEUM|MESOTHELIOMA OF MESOCOLON
C0496767|T191|C10.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF OROPHARYNX|BOESARTIGE NEUBILDUNG: OROPHARYNX, MEHRERE TEILBEREICHE UEBERLAPPEND
C0153382|T191|C10.9|DMDICD10|MALIGNANT NEOPLASM OF OROPHARYNX, UNSPECIFIED|BOESARTIGE NEUBILDUNG: OROPHARYNX, NICHT NAEHER BEZEICHNET
C2833847|T191|C10.4|ICD10CM|MALIGNANT NEOPLASM OF BRANCHIAL CLEFT|MALIGNANT NEOPLASM OF BRANCHIAL CYST [SITE OF NEOPLASM]
C0025500|T191|C45.9|DMDICD10|MESOTHELIOMA, UNSPECIFIED|MESOTHELIOM, NICHT NAEHER BEZEICHNET
C0153386|T191|C10.0|DMDICD10|MALIGNANT NEOPLASM OF VALLECULA|BOESARTIGE NEUBILDUNG: VALLECULA EPIGLOTTICA
C2833846|T191|C10.1|ICD10CM|MALIGNANT NEOPLASM OF ANTERIOR SURFACE OF EPIGLOTTIS|MALIGNANT NEOPLASM OF EPIGLOTTIS, FREE BORDER [MARGIN]
C0153389|T191|C10.2|DMDICD10|MALIGNANT NEOPLASM OF LATERAL WALL OF OROPHARYNX|BOESARTIGE NEUBILDUNG: SEITENWAND DES OROPHARYNX
C0153390|T191|C10.3|DMDICD10|MALIGNANT NEOPLASM OF POSTERIOR WALL OF OROPHARYNX|BOESARTIGE NEUBILDUNG: HINTERWAND DES OROPHARYNX
C2861677|T191|D03.60|ICD10CM|MELANOMA IN SITU OF UNSPECIFIED UPPER LIMB, INCLUDING SHOULDER|MELANOMA IN SITU OF UNSP UPPER LIMB, INCLUDING SHOULDER
C2861678|T191|D03.61|ICD10CM|MELANOMA IN SITU OF RIGHT UPPER LIMB, INCLUDING SHOULDER|MELANOMA IN SITU OF RIGHT UPPER LIMB, INCLUDING SHOULDER
C2861679|T191|D03.62|ICD10CM|MELANOMA IN SITU OF LEFT UPPER LIMB, INCLUDING SHOULDER|MELANOMA IN SITU OF LEFT UPPER LIMB, INCLUDING SHOULDER
C2874494|T048|F12.280|ICD10CM|CANNABIS DEPENDENCE WITH CANNABIS-INDUCED ANXIETY DISORDER|CANNABIS DEPENDENCE WITH CANNABIS-INDUCED ANXIETY DISORDER
C2832313|T037|S06.362A|ICD10CM|TRAUMATIC HEMORRHAGE OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|TRAUM HEMOR CEREB, W LOC OF 31-59 MIN, INIT
C2890809|T037|T84.52XA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL LEFT HIP PROSTHESIS, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INTERNAL LEFT HIP PROSTH, INIT
C2890555|T037|T84.090A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTERNAL RIGHT HIP PROSTHESIS, INITIAL ENCOUNTER|MECH COMPL OF INTERNAL RIGHT HIP PROSTHESIS, INIT ENCNTR
C2832315|T037|S06.362S|ICD10CM|TRAUMATIC HEMORRHAGE OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|TRAUM HEMOR CEREB, W LOC OF 31-59 MIN, SEQUELA
C0348469|T047|E22|DMDICD10|HYPERFUNCTION OF PITUITARY GLAND, UNSPECIFIED|UEBERFUNKTION DER HYPOPHYSE
C0348456|T046|E22.8|DMDICD10|OTHER HYPERFUNCTION OF PITUITARY GLAND|SONSTIGE UEBERFUNKTION DER HYPOPHYSE
C2832115|T037|S06.315A|ICD10CM|CONTUSION AND LACERATION OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, INITIAL ENCOUNTER|CONTUS/LAC RIGHT CEREBRUM W LOC >24 HR W RET CONSC LEV, INIT
C2857564|T037|S72.21XA|ICD10CM|DISPLACED SUBTROCHANTERIC FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED SUBTROCHANTERIC FRACTURE OF RIGHT FEMUR, INIT
C0021141|T047|E22.2|DMDICD10|SYNDROME OF INAPPROPRIATE SECRETION OF ANTIDIURETIC HORMONE|SYNDROM DER INADAEQUATEN SEKRETION VON ADIURETIN
C0020514|T047|E22.1|DMDICD10|HYPERPROLACTINEMIA|HYPERPROLAKTINAEMIE
C0405578|T047|E22.0|DMDICD10|ACROMEGALY AND PITUITARY GIGANTISM|AKROMEGALIE UND HYPOPHYSAERER RIESENWUCHS
C2838257|T037|S32.466A|ICD10CM|NONDISPLACED ASSOCIATED TRANSVERSE-POSTERIOR FRACTURE OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP ASSOCIATED TRANSV/POST FX UNSP ACETABULUM, INIT
C2857566|T037|S72.21XC|ICD10CM|DISPLACED SUBTROCHANTERIC FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPLACED SUBTROCHNT FX R FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C1455979|T033|Z79.4|ICD10CM|LONG TERM (CURRENT) USE OF INSULIN|LONG TERM (CURRENT) USE OF INSULIN
C2832356|T037|S06.372S|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF CEREBELLUM WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|CONTUS/LAC/HEM CRBLM W LOC OF 31-59 MIN, SEQUELA
C2977643|T033|Z68.41|ICD10CM|BODY MASS INDEX (BMI) 40.0-44.9, ADULT|BODY MASS INDEX (BMI) 40.0-44.9, ADULT
C2887912|T047|K70.30|ICD10CM|ALCOHOLIC CIRRHOSIS OF LIVER WITHOUT ASCITES|ALCOHOLIC CIRRHOSIS OF LIVER WITHOUT ASCITES
C2887913|T047|K70.31|ICD10CM|ALCOHOLIC CIRRHOSIS OF LIVER WITH ASCITES|ALCOHOLIC CIRRHOSIS OF LIVER WITH ASCITES
C2832354|T037|S06.372A|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF CEREBELLUM WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|CONTUS/LAC/HEM CRBLM W LOC OF 31-59 MIN, INIT
C4270383|T046|T83.714A|ICD10CM|EROSION OF IMPLANTED URETERAL BULKING AGENT TO SURROUNDING ORGAN OR TISSUE, INITIAL ENCOUNTER|EROSN IMPLNT URTL BULK AGNT ORGAN OR TISSUE, INIT
C2977646|T033|Z68.44|ICD10CM|BODY MASS INDEX (BMI) 60.0-69.9, ADULT|BODY MASS INDEX (BMI) 60.0-69.9, ADULT
C2888352|T047|L89.153|ICD10CM|PRESSURE ULCER OF SACRAL REGION, STAGE 3|PRESSURE ULCER OF SACRAL REGION, STAGE 3
C2888349|T047|L89.152|ICD10CM|PRESSURE ULCER OF SACRAL REGION, STAGE 2|PRESSURE ULCER OF SACRAL REGION, STAGE 2
C2888346|T047|L89.151|ICD10CM|PRESSURE ULCER OF SACRAL REGION, STAGE 1|PRESSURE ULCER OF SACRAL REGION, STAGE 1
C2888343|T047|L89.150|ICD10CM|PRESSURE ULCER OF SACRAL REGION, UNSTAGEABLE|PRESSURE ULCER OF SACRAL REGION, UNSTAGEABLE
C2888355|T047|L89.154|ICD10CM|PRESSURE ULCER OF SACRAL REGION, STAGE 4|PRESSURE ULCER OF SACRAL REGION, STAGE 4
C2861624|T191||ICD10CM|JUVENILE MYELOMONOCYTIC LEUKEMIA, IN RELAPSE
C2888358|T047|L89.159|ICD10CM|PRESSURE ULCER OF SACRAL REGION, UNSPECIFIED STAGE|PRESSURE ULCER OF SACRAL REGION, UNSPECIFIED STAGE
C2861622|T191|C93.30|ICD10CM|JUVENILE MYELOMONOCYTIC LEUKEMIA, NOT HAVING ACHIEVED REMISSION|JUVENILE MYELOMONOCYTIC LEUKEMIA, NOT ACHIEVE REMISSION
C2837869|T037|S32.391B|ICD10CM|OTHER FRACTURE OF RIGHT ILIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTHER FRACTURE OF RIGHT ILIUM, INIT ENCNTR FOR OPEN FRACTURE
C0339963|T047|B38.1|DMDICD10|CHRONIC PULMONARY COCCIDIOIDOMYCOSIS|CHRONISCHE KOKZIDIOIDOMYKOSE DER LUNGE
C2882493|T047|I69.131|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING RIGHT DOMINANT SIDE|MONOPLG UPR LMB FOL NTRM INTCRBL HEMOR AFF RIGHT DOM SIDE
C2882494|T047|I69.132|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING LEFT DOMINANT SIDE|MONOPLG UPR LMB FOL NTRM INTCRBL HEMOR AFF LEFT DOM SIDE
C0375046|T047|B38.2|DMDICD10|PULMONARY COCCIDIOIDOMYCOSIS, UNSPECIFIED|KOKZIDIOIDOMYKOSE DER LUNGE, NICHT NAEHER BEZEICHNET
C2889471|T047|M06.821|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, RIGHT ELBOW|OTHER SPECIFIED RHEUMATOID ARTHRITIS, RIGHT ELBOW
C2902431|T047|M90.529|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, UNSPECIFIED UPPER ARM|OSTEONECROSIS IN DISEASES CLASSD ELSWHR, UNSP UPPER ARM
C2889472|T047|M06.822|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, LEFT ELBOW|OTHER SPECIFIED RHEUMATOID ARTHRITIS, LEFT ELBOW
C2882497|T047|I69.139|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING UNSPECIFIED SIDE|MONOPLG UPR LMB FOLLOWING NTRM INTCRBL HEMOR AFF UNSP SIDE
C2889473|T047|M06.829|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, UNSPECIFIED ELBOW|OTHER SPECIFIED RHEUMATOID ARTHRITIS, UNSPECIFIED ELBOW
C2874836|T048|F19.920|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH INTOXICATION, UNCOMPLICATED|OTH PSYCHOACTIVE SUBSTANCE USE, UNSP W INTOXICATION, UNCOMP
C2902429|T047|M90.521|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, RIGHT UPPER ARM|OSTEONECROSIS IN DISEASES CLASSD ELSWHR, RIGHT UPPER ARM
C2874838|T048|F19.922|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE|OTH PSYCHOACTV SUB USE, UNSP W INTOX W PERCEPTL DISTURB
C2886033|T037|T65.222A|ICD10CM|TOXIC EFFECT OF TOBACCO CIGARETTES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF TOBACCO CIGARETTES, SELF-HARM, INIT
C2889606|T047|M08.829|ICD10CM|OTHER JUVENILE ARTHRITIS, UNSPECIFIED ELBOW|OTHER JUVENILE ARTHRITIS, UNSPECIFIED ELBOW
C2857377|T037|S72.132A|ICD10CM|DISPLACED APOPHYSEAL FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED APOPHYSEAL FRACTURE OF LEFT FEMUR, INIT
C2889605|T047|M08.822|ICD10CM|OTHER JUVENILE ARTHRITIS, LEFT ELBOW|OTHER JUVENILE ARTHRITIS, LEFT ELBOW
C2889604|T047|M08.821|ICD10CM|OTHER JUVENILE ARTHRITIS, RIGHT ELBOW|OTHER JUVENILE ARTHRITIS, RIGHT ELBOW
C2857378|T037|S72.132B|ICD10CM|DISPLACED APOPHYSEAL FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPLACED APOPHYSEAL FX LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C0349368|T047|I15.2|DMDICD10|HYPERTENSION SECONDARY TO ENDOCRINE DISORDERS|HYPERTONIE ALS FOLGE VON ENDOKRINEN KRANKHEITEN
C2901911|T047|M86.572|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, LEFT ANKLE AND FOOT|OTH CHRONIC HEMATOGENOUS OSTEOMYELITIS, LEFT ANKLE AND FOOT
C2901910|T047|M86.571|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, RIGHT ANKLE AND FOOT|OTH CHRONIC HEMATOGENOUS OSTEOMYELITIS, RIGHT ANKLE AND FOOT
C2901912|T047|M86.579|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED ANKLE AND FOOT|OTH CHRONIC HEMATOGENOUS OSTEOMYELITIS, UNSP ANKLE AND FOOT
C2885475|T037|T63.122A|ICD10CM|TOXIC EFFECT OF VENOM OF OTHER VENOMOUS LIZARD, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF VENOMOUS LIZARD, SELF-HARM, INIT
C2885477|T037|T63.122S|ICD10CM|TOXIC EFFECT OF VENOM OF OTHER VENOMOUS LIZARD, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF VENOMOUS LIZARD, SELF-HARM, SEQUELA
C2833777|T037|S14.101S|ICD10CM|UNSPECIFIED INJURY AT C1 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|UNSP INJURY AT C1 LEVEL OF CERVICAL SPINAL CORD, SEQUELA
C2877591|T037|T40.1X2S|ICD10CM|POISONING BY HEROIN, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY HEROIN, INTENTIONAL SELF-HARM, SEQUELA
C2877613|T037|T40.2X2A|ICD10CM|POISONING BY OTHER OPIOIDS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH OPIOIDS, INTENTIONAL SELF-HARM, INIT ENCNTR
C2833775|T037|S14.101A|ICD10CM|UNSPECIFIED INJURY AT C1 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY AT C1 LEVEL OF CERVICAL SPINAL CORD, INIT ENCNTR
C2865589|T037|S88.929A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED LOWER LEG, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP OF UNSP LOWER LEG, LEVEL UNSP, INIT
C2877615|T037|T40.2X2S|ICD10CM|POISONING BY OTHER OPIOIDS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTHER OPIOIDS, INTENTIONAL SELF-HARM, SEQUELA
C2833776|T037|S14.101D|ICD10CM|UNSPECIFIED INJURY AT C1 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY AT C1 LEVEL OF CERVICAL SPINAL CORD, SUBS ENCNTR
C2242472|T047||ICD10CM|OSTEOMYELITIS, UNSPECIFIED
C2858976|T037|S72.491A|ICD10CM|OTHER FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF LOWER END OF RIGHT FEMUR, INIT FOR CLOS FX
C2885356|T037|T63.032A|ICD10CM|TOXIC EFFECT OF TAIPAN VENOM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF TAIPAN VENOM, INTENTIONAL SELF-HARM, INIT
C2858978|T037|S72.491C|ICD10CM|OTHER FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|OTH FX LOWER END OF RIGHT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2858977|T037|S72.491B|ICD10CM|OTHER FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|OTH FX LOWER END OF RIGHT FEMUR, INIT FOR OPN FX TYPE I/2
C2858406|T037|S72.415A|ICD10CM|NONDISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP UNSP CONDYLE FX LOWER END OF LEFT FEMUR, INIT
C3264226|T047|H40.1390|ICD10CM|PIGMENTARY GLAUCOMA, UNSPECIFIED EYE, STAGE UNSPECIFIED|PIGMENTARY GLAUCOMA, UNSPECIFIED EYE, STAGE UNSPECIFIED
C3264227|T047|H40.1391|ICD10CM|PIGMENTARY GLAUCOMA, UNSPECIFIED EYE, MILD STAGE|PIGMENTARY GLAUCOMA, UNSPECIFIED EYE, MILD STAGE
C3264228|T047|H40.1392|ICD10CM|PIGMENTARY GLAUCOMA, UNSPECIFIED EYE, MODERATE STAGE|PIGMENTARY GLAUCOMA, UNSPECIFIED EYE, MODERATE STAGE
C3264229|T047|H40.1393|ICD10CM|PIGMENTARY GLAUCOMA, UNSPECIFIED EYE, SEVERE STAGE|PIGMENTARY GLAUCOMA, UNSPECIFIED EYE, SEVERE STAGE
C3264230|T047|H40.1394|ICD10CM|PIGMENTARY GLAUCOMA, UNSPECIFIED EYE, INDETERMINATE STAGE|PIGMENTARY GLAUCOMA, UNSPECIFIED EYE, INDETERMINATE STAGE
C2865585|T037|S88.922A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT LOWER LEG, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF L LOW LEG, LEVEL UNSP, INIT
C2865586|T037|S88.922D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT LOWER LEG, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF L LOW LEG, LEVEL UNSP, SUBS
C2832531|T037|S06.6X5S|ICD10CM|TRAUMATIC SUBARACHNOID HEMORRHAGE WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, SEQUELA|TRAUM SUBRAC HEM W LOC >24 HR W RET CONSC LEV, SEQUELA
C2865587|T037|S88.922S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT LOWER LEG, LEVEL UNSPECIFIED, SEQUELA|PARTIAL TRAUMATIC AMP OF L LOW LEG, LEVEL UNSP, SEQUELA
C2880024|T037|T48.3X2A|ICD10CM|POISONING BY ANTITUSSIVES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ANTITUSSIVES, INTENTIONAL SELF-HARM, INIT
C2832529|T037|S06.6X5A|ICD10CM|TRAUMATIC SUBARACHNOID HEMORRHAGE WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, INITIAL ENCOUNTER|TRAUM SUBRAC HEM W LOC >24 HR W RET CONSC LEV, INIT
C0086795|T047||ICD10CM|HURLER'S SYNDROME
C2838086|T037|S32.426B|ICD10CM|NONDISPLACED FRACTURE OF POSTERIOR WALL OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP FX OF POSTERIOR WALL OF UNSP ACETAB, INIT FOR OPN FX
C4268408|T047|H40.1134|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, BILATERAL, INDETERMINATE STAGE|PRIMARY OPEN-ANGLE GLAUCOMA, BILATERAL, INDETERMINATE STAGE
C2889172|T047|M05.229|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF UNSP ELBOW
C4268404|T047|H40.1130|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, BILATERAL, STAGE UNSPECIFIED|PRIMARY OPEN-ANGLE GLAUCOMA, BILATERAL, STAGE UNSPECIFIED
C4268405|T047|H40.1131|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, BILATERAL, MILD STAGE|PRIMARY OPEN-ANGLE GLAUCOMA, BILATERAL, MILD STAGE
C4268406|T047|H40.1132|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, BILATERAL, MODERATE STAGE|PRIMARY OPEN-ANGLE GLAUCOMA, BILATERAL, MODERATE STAGE
C4268407|T047|H40.1133|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, BILATERAL, SEVERE STAGE|PRIMARY OPEN-ANGLE GLAUCOMA, BILATERAL, SEVERE STAGE
C2882770|T047|I70.334|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF HEEL AND MIDFOOT|ATHSCL UNSP TYPE BYPASS OF R LEG W ULCER OF HEEL AND MIDFT
C2882772|T047|I70.335|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF OTHER PART OF FOOT|ATHSCL UNSP TYPE BYPASS OF RIGHT LEG W ULCER OTH PRT FOOT
C2889170|T047|M05.221|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT ELBOW|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF RIGHT ELBOW
C2905705|T037|X74.02XS|ICD10CM|INTENTIONAL SELF-HARM BY PAINTBALL GUN, SEQUELA|INTENTIONAL SELF-HARM BY PAINTBALL GUN, SEQUELA
C2882766|T047|I70.331|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF THIGH|ATHSCL UNSP TYPE BYPASS OF THE RIGHT LEG W ULCER OF THIGH
C2882767|T047|I70.332|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF CALF|ATHSCL UNSP TYPE BYPASS OF THE RIGHT LEG W ULCER OF CALF
C2882768|T047|I70.333|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF ANKLE|ATHSCL UNSP TYPE BYPASS OF THE RIGHT LEG W ULCER OF ANKLE
C2865542|T037|S88.111A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, RIGHT LOWER LEG, INITIAL ENCOUNTER|COMPLETE TRAUM AMP AT LEV BETW KN AND ANKL, R LOW LEG, INIT
C2905734|T037|X77.2XXA|ICD10CM|INTENTIONAL SELF-HARM BY OTHER HOT FLUIDS, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY OTHER HOT FLUIDS, INITIAL ENCOUNTER
C2865543|T037|S88.111D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, RIGHT LOWER LEG, SUBSEQUENT ENCOUNTER|COMPLETE TRAUM AMP AT LEV BETW KN AND ANKL, R LOW LEG, SUBS
C2905735|T037|X77.2XXD|ICD10CM|INTENTIONAL SELF-HARM BY OTHER HOT FLUIDS, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY OTHER HOT FLUIDS, SUBS ENCNTR
C2832645|T037|S06.893S|ICD10CM|OTHER SPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, SEQUELA|INTCRAN INJ W LOC OF 1-5 HRS 59 MIN, SEQUELA
C2500065|T060|B20|ICD10PCS|HUMAN IMMUNODEFICIENCY VIRUS [HIV] DISEASE|IMAGING @ HEART @ PLAIN RADIOGRAPHY
C2905736|T037|X77.2XXS|ICD10CM|INTENTIONAL SELF-HARM BY OTHER HOT FLUIDS, SEQUELA|INTENTIONAL SELF-HARM BY OTHER HOT FLUIDS, SEQUELA
C2865544|T037|S88.111S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, RIGHT LOWER LEG, SEQUELA|COMPLETE TRAUM AMP AT LEV BETW KN AND ANKL, R LOW LEG, SQLA
C0242770|T047||ICD10CM|CRYPTOGENIC ORGANIZING PNEUMONIA
C0238378|T047|J84.117|ICD10CM|DESQUAMATIVE INTERSTITIAL PNEUMONIA|DESQUAMATIVE INTERSTITIAL PNEUMONIA
C1279945|T047|J84.114|ICD10CM|ACUTE INTERSTITIAL PNEUMONITIS|ACUTE INTERSTITIAL PNEUMONITIS
C0238378|T047|J84.117|ICD10CM|RESPIRATORY BRONCHIOLITIS INTERSTITIAL LUNG DISEASE|DESQUAMATIVE INTERSTITIAL PNEUMONIA
C1800706|T047||ICD10CM|IDIOPATHIC PULMONARY FIBROSIS
C3161102|T047|J84.113|ICD10CM|IDIOPATHIC NON-SPECIFIC INTERSTITIAL PNEUMONITIS|IDIOPATHIC NON-SPECIFIC INTERSTITIAL PNEUMONITIS
C4270379|T046|T83.713A|ICD10CM|EROSION OF IMPLANTED URETHRAL BULKING AGENT TO SURROUNDING ORGAN OR TISSUE, INITIAL ENCOUNTER|EROSN IMPLNT URETHRAL BULKING AGENT TO SURRND ORG/TISS, INIT
C3161100|T046|J84.111|ICD10CM|IDIOPATHIC INTERSTITIAL PNEUMONIA, NOT OTHERWISE SPECIFIED|IDIOPATHIC INTERSTITIAL PNEUMONIA, NOT OTHERWISE SPECIFIED
C2884002|T037|T51.1X2A|ICD10CM|TOXIC EFFECT OF METHANOL, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF METHANOL, INTENTIONAL SELF-HARM, INIT ENCNTR
C2869870|T037|S98.319D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED MIDFOOT, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF UNSP MIDFOOT, SUBS ENCNTR
C2869869|T037|S98.319A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED MIDFOOT, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF UNSP MIDFOOT, INIT ENCNTR
C2838366|T037|S32.499B|ICD10CM|OTHER SPECIFIED FRACTURE OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF UNSP ACETABULUM, INIT FOR OPN FX
C2845896|T191|C66.1|ICD10CM|MALIGNANT NEOPLASM OF RIGHT URETER|MALIGNANT NEOPLASM OF RIGHT URETER
C2858937|T037|S72.466B|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP SUPRCNDL FX W INTRCNDL EXTN LOW END UNSP FEMR, 7THB
C2858936|T037|S72.466A|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP SUPRCNDL FX W INTRCNDL EXTN LOW END UNSP FEMR, INIT
C2977943|T191|C66.2|ICD10CM|MALIGNANT NEOPLASM OF LEFT URETER|MALIGNANT NEOPLASM OF LEFT URETER
C2902430|T047|M90.522|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, LEFT UPPER ARM|OSTEONECROSIS IN DISEASES CLASSD ELSWHR, LEFT UPPER ARM
C2845897|T191|C66.9|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED URETER|MALIGNANT NEOPLASM OF UNSPECIFIED URETER
C2902739|T037|M96.669|ICD10CM|FRACTURE OF FEMUR FOLLOWING INSERTION OF ORTHOPEDIC IMPLANT, JOINT PROSTHESIS, OR BONE PLATE, UNSPECIFIED LEG|FX FEMUR FOL INSRT ORTHO IMPLNT/PROSTH/BONE PLT, UNSP LEG
C0023788|T047||ICD10CM|WHIPPLE'S DISEASE
C2885886|T037|T63.822S|ICD10CM|TOXIC EFFECT OF CONTACT WITH VENOMOUS TOAD, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CONTACT W VENOMOUS TOAD, SELF-HARM, SEQUELA
C0341288|T047|K90.8|ICD10CM|OTHER INTESTINAL MALABSORPTION|OTHER INTESTINAL MALABSORPTION
C2838158|T037|S32.444B|ICD10CM|NONDISPLACED FRACTURE OF POSTERIOR COLUMN [ILIOISCHIAL] OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP FX OF POST COLUMN OF RIGHT ACETAB, INIT FOR OPN FX
C0494273|T047|E03.8|DMDICD10|OTHER SPECIFIED HYPOTHYROIDISM|SONSTIGE NAEHER BEZEICHNETE HYPOTHYREOSE
C0027145|T047||ICD10CM|HYPOTHYROIDISM, UNSPECIFIED
C0342197|T020|E03.4|DMDICD10|ATROPHY OF THYROID (ACQUIRED)|ATROPHIE DER SCHILDDRUESE (ERWORBEN)
C0238298|T047|E03.5|DMDICD10|MYXEDEMA COMA|MYXOEDEMKOMA
C0494272|T047|E03.2|DMDICD10|HYPOTHYROIDISM DUE TO MEDICAMENTS AND OTHER EXOGENOUS SUBSTANCES|HYPOTHYREOSE DURCH ARZNEIMITTEL ODER ANDERE EXOGENE SUBSTANZEN
C0342173|T047|E03.3|DMDICD10|POSTINFECTIOUS HYPOTHYROIDISM|POSTINFEKTIOESE HYPOTHYREOSE
C2873860|T046|E03.0|ICD10CM|CONGENITAL HYPOTHYROIDISM WITH DIFFUSE GOITER|CONGENITAL PARENCHYMATOUS GOITER (NONTOXIC)
C0749420|T019||ICD10CM|CONGENITAL HYPOTHYROIDISM WITHOUT GOITER
C2874196|T047|E27.49|ICD10CM|OTHER ADRENOCORTICAL INSUFFICIENCY|OTHER ADRENOCORTICAL INSUFFICIENCY
C0020595|T047|E27.40|ICD10CM|UNSPECIFIED ADRENOCORTICAL INSUFFICIENCY|UNSPECIFIED ADRENOCORTICAL INSUFFICIENCY
C2874636|T048|F15.15|ICD10CM|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER
C2857771|T037|S72.324B|ICD10CM|NONDISPLACED TRANSVERSE FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP TRANSVERSE FX SHAFT OF R FEMR, 7THB
C2857772|T037|S72.324C|ICD10CM|NONDISPLACED TRANSVERSE FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP TRANSVERSE FX SHAFT OF R FEMR, 7THC
C2833479|T037|S12.44XA|ICD10CM|TYPE III TRAUMATIC SPONDYLOLISTHESIS OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE III TRAUM SPONDYLOLYSIS OF FIFTH CERVCAL VERTEBRA, INIT
C2586056|T046|I48.2|ICD10CM|CHRONIC ATRIAL FIBRILLATION|PERMANENT ATRIAL FIBRILLATION
C2874634|T048|F15.150|ICD10CM|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|OTH STIMULANT ABUSE W STIM-INDUCE PSYCH DISORDER W DELUSIONS
C2874635|T048|F15.151|ICD10CM|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|OTH STIMULANT ABUSE W STIM-INDUCE PSYCH DISORDER W HALLUCIN
C2585653|T046|I48.1|ICD10CM|PERSISTENT ATRIAL FIBRILLATION|PERSISTENT ATRIAL FIBRILLATION
C2845969|T191|C79.40|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF UNSPECIFIED PART OF NERVOUS SYSTEM|SECONDARY MALIGNANT NEOPLASM OF UNSP PART OF NERVOUS SYSTEM
C2875366|T047|G90.3|ICD10CM|MULTI-SYSTEM DEGENERATION OF THE AUTONOMIC NERVOUS SYSTEM|MULTI-SYSTEM DEGENERATION OF THE AUTONOMIC NERVOUS SYSTEM
C2877815|T037|T40.902A|ICD10CM|POISONING BY UNSPECIFIED PSYCHODYSLEPTICS [HALLUCINOGENS], INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY UNSP PSYCHODYSLEPTICS, SELF-HARM, INIT
C2890300|T037|T83.22XA|ICD10CM|DISPLACEMENT OF GRAFT OF URINARY ORGAN, INITIAL ENCOUNTER|DISPLACEMENT OF GRAFT OF URINARY ORGAN, INITIAL ENCOUNTER
C0153689|T191|C79.49|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF OTHER PARTS OF NERVOUS SYSTEM|SECONDARY MALIGNANT NEOPLASM OF OTH PARTS OF NERVOUS SYSTEM
C2895311|T037|M48.50XA|ICD10CM|COLLAPSED VERTEBRA, NOT ELSEWHERE CLASSIFIED, SITE UNSPECIFIED, INITIAL ENCOUNTER FOR FRACTURE|COLLAPSED VERTEBRA, NEC, SITE UNSP, INIT
C2910018|T047|P36.19|ICD10CM|SEPSIS OF NEWBORN DUE TO OTHER STREPTOCOCCI|SEPSIS OF NEWBORN DUE TO OTHER STREPTOCOCCI
C2877817|T037|T40.902S|ICD10CM|POISONING BY UNSPECIFIED PSYCHODYSLEPTICS [HALLUCINOGENS], INTENTIONAL SELF-HARM, SEQUELA|POISONING BY UNSP PSYCHODYSLEPTICS, SELF-HARM, SEQUELA
C2830350|T033|R40.2111|ICD10CM|COMA SCALE, EYES OPEN, NEVER, IN THE FIELD [EMT OR AMBULANCE]|COMA SCALE, EYES OPEN, NEVER, IN THE FIELD
C2830349|T033|R40.2110|ICD10CM|COMA SCALE, EYES OPEN, NEVER, UNSPECIFIED TIME|COMA SCALE, EYES OPEN, NEVER, UNSPECIFIED TIME
C2830352|T033|R40.2113|ICD10CM|COMA SCALE, EYES OPEN, NEVER, AT HOSPITAL ADMISSION|COMA SCALE, EYES OPEN, NEVER, AT HOSPITAL ADMISSION
C2830351|T033|R40.2112|ICD10CM|COMA SCALE, EYES OPEN, NEVER, AT ARRIVAL TO EMERGENCY DEPARTMENT|COMA SCALE, EYES OPEN, NEVER, EMR
C2830353|T033|R40.2114|ICD10CM|COMA SCALE, EYES OPEN, NEVER, 24 HOURS OR MORE AFTER HOSPITAL ADMISSION|COMA SCALE, EYES OPEN, NEVER, 24+HRS
C2883535|T037|T50.0X2S|ICD10CM|POISONING BY MINERALOCORTICOIDS AND THEIR ANTAGONISTS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY MINERALOCORTICOIDS AND ANTAG, SELF-HARM, SEQUELA
C0154120|T191|D42.9|DMDICD10|NEOPLASM OF UNCERTAIN BEHAVIOR OF MENINGES, UNSPECIFIED|NEUBILDUNG UNSICHEREN ODER UNBEKANNTEN VERHALTENS: MENINGEN, NICHT NAEHER BEZEICHNET
C2838502|T037|S32.811A|ICD10CM|MULTIPLE FRACTURES OF PELVIS WITH UNSTABLE DISRUPTION OF PELVIC RING, INITIAL ENCOUNTER FOR CLOSED FRACTURE|MULT FX OF PELVIS W UNSTABLE DISRUPT OF PELVIC RING, INIT
C2838503|T037|S32.811B|ICD10CM|MULTIPLE FRACTURES OF PELVIS WITH UNSTABLE DISRUPTION OF PELVIC RING, INITIAL ENCOUNTER FOR OPEN FRACTURE|MULT FX OF PELV W UNSTBL DISRUPT OF PELV RING, 7THB
C2838458|T037|S32.615B|ICD10CM|NONDISPLACED AVULSION FRACTURE OF LEFT ISCHIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP AVULSION FRACTURE OF LEFT ISCHIUM, INIT FOR OPN FX
C2838457|T037|S32.615A|ICD10CM|NONDISPLACED AVULSION FRACTURE OF LEFT ISCHIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED AVULSION FRACTURE OF LEFT ISCHIUM, INIT
C2869834|T037|S98.211A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF TWO OR MORE RIGHT LESSER TOES, INITIAL ENCOUNTER|COMPLETE TRAUM AMP OF TWO OR MORE RIGHT LESSER TOES, INIT
C1719322|T047|D61.09|ICD10CM|OTHER CONSTITUTIONAL APLASTIC ANEMIA|OTHER CONSTITUTIONAL APLASTIC ANEMIA
C2869835|T037|S98.211D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF TWO OR MORE RIGHT LESSER TOES, SUBSEQUENT ENCOUNTER|COMPLETE TRAUM AMP OF TWO OR MORE RIGHT LESSER TOES, SUBS
C2874115|T047|E11.621|ICD10CM|TYPE 2 DIABETES MELLITUS WITH FOOT ULCER|TYPE 2 DIABETES MELLITUS WITH FOOT ULCER
C2869836|T037|S98.211S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF TWO OR MORE RIGHT LESSER TOES, SEQUELA|COMPLETE TRAUM AMP OF TWO OR MORE RIGHT LESSER TOES, SEQUELA
C2874114|T047|E11.620|ICD10CM|TYPE 2 DIABETES MELLITUS WITH DIABETIC DERMATITIS|TYPE 2 DIABETES MELLITUS WITH DIABETIC DERMATITIS
C2856045|T037|S68.620S|ICD10CM|PARTIAL TRAUMATIC TRANSPHALANGEAL AMPUTATION OF RIGHT INDEX FINGER, SEQUELA|PARTIAL TRAUMATIC TRNSPHAL AMPUTATION OF R IDX FNGR, SEQUELA
C2848417|T037|S58.111S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN ELBOW AND WRIST, RIGHT ARM, SEQUELA|COMPLETE TRAUM AMP AT LEV BETW ELBOW AND WRIST, R ARM, SQLA
C2905664|T037|X71.8XXS|ICD10CM|OTHER INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION, SEQUELA|OTH INTENTIONAL SELF-HARM BY DROWN, SEQUELA
C2888528|T047|L89.529|ICD10CM|PRESSURE ULCER OF LEFT ANKLE, UNSPECIFIED STAGE|PRESSURE ULCER OF LEFT ANKLE, UNSPECIFIED STAGE
C2888519|T047|L89.522|ICD10CM|PRESSURE ULCER OF LEFT ANKLE, STAGE 2|PRESSURE ULCER OF LEFT ANKLE, STAGE 2
C2888522|T047|L89.523|ICD10CM|PRESSURE ULCER OF LEFT ANKLE, STAGE 3|PRESSURE ULCER OF LEFT ANKLE, STAGE 3
C2888513|T047||ICD10CM|PRESSURE ULCER OF LEFT ANKLE, UNSTAGEABLE
C4268683|T047|L89.521|ICD10CM|PRESSURE ULCER OF LEFT ANKLE, STAGE 1|PRESSURE PRE-ULCER SKIN CHANGES LIMITED TO PERSISTENT FOCAL EDEMA, LEFT ANKLE
C2888525|T047|L89.524|ICD10CM|PRESSURE ULCER OF LEFT ANKLE, STAGE 4|PRESSURE ULCER OF LEFT ANKLE, STAGE 4
C2882968|T047|I70.693|ICD10CM|OTHER ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, BILATERAL LEGS|OTH ATHSCL NONBIOL BYPASS OF THE EXTREMITIES, BILATERAL LEGS
C2882967|T047|I70.692|ICD10CM|OTHER ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, LEFT LEG|OTH ATHSCL NONBIOLOGICAL BYPASS OF THE EXTREMITIES, LEFT LEG
C2882966|T047|I70.691|ICD10CM|OTHER ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, RIGHT LEG|OTH ATHSCL NONBIOL BYPASS OF THE EXTREMITIES, RIGHT LEG
C2874687|T048|F16.151|ICD10CM|HALLUCINOGEN ABUSE WITH HALLUCINOGEN-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|HALLUCINOGEN ABUSE W PSYCHOTIC DISORDER W HALLUCINATIONS
C2874686|T048|F16.150|ICD10CM|HALLUCINOGEN ABUSE WITH HALLUCINOGEN-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|HALLUCINOGEN ABUSE W PSYCHOTIC DISORDER W DELUSIONS
C0838502|T047|M46.20|ICD10AM|OSTEOMYELITIS OF VERTEBRA, SITE UNSPECIFIED|OSTEOMYELITIS OF VERTEBRA, MULTIPLE SITES IN SPINE
C0838503|T047|M46.21|ICD10AM|OSTEOMYELITIS OF VERTEBRA, OCCIPITO-ATLANTO-AXIAL REGION|OSTEOMYELITIS OF VERTEBRA, OCCIPITO-ATLANTO-AXIAL REGION
C2882970|T047|I70.699|ICD10CM|OTHER ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, UNSPECIFIED EXTREMITY|OTH ATHSCL NONBIOL BYPASS OF THE EXTREMITIES, UNSP EXTREMITY
C2882969|T047|I70.698|ICD10CM|OTHER ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, OTHER EXTREMITY|OTH ATHSCL NONBIOL BYPASS OF THE EXTREMITIES, OTH EXTREMITY
C2874688|T048|F16.159|ICD10CM|HALLUCINOGEN ABUSE WITH HALLUCINOGEN-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|HALLUCINOGEN ABUSE WITH HALLUCINOGEN-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED
C0838507|T047|M46.25|ICD10AM|OSTEOMYELITIS OF VERTEBRA, THORACOLUMBAR REGION|OSTEOMYELITIS OF VERTEBRA, THORACOLUMBAR REGION
C0838508|T047|M46.26|ICD10AM|OSTEOMYELITIS OF VERTEBRA, LUMBAR REGION|OSTEOMYELITIS OF VERTEBRA, LUMBAR REGION
C0838509|T047|M46.27|ICD10AM|OSTEOMYELITIS OF VERTEBRA, LUMBOSACRAL REGION|OSTEOMYELITIS OF VERTEBRA, LUMBOSACRAL REGION
C0348457|T047|E23.6|DMDICD10|OTHER DISORDERS OF PITUITARY GLAND|SONSTIGE STOERUNGEN DER HYPOPHYSE
C2888850|T047|M00.162|ICD10CM|PNEUMOCOCCAL ARTHRITIS, LEFT KNEE|PNEUMOCOCCAL ARTHRITIS, LEFT KNEE
C2874050|T047|E10.49|ICD10CM|TYPE 1 DIABETES MELLITUS WITH OTHER DIABETIC NEUROLOGICAL COMPLICATION|TYPE 1 DIABETES W OTH DIABETIC NEUROLOGICAL COMPLICATION
C2888849|T047|M00.161|ICD10CM|PNEUMOCOCCAL ARTHRITIS, RIGHT KNEE|PNEUMOCOCCAL ARTHRITIS, RIGHT KNEE
C2874048|T047|E10.43|ICD10CM|TYPE 1 DIABETES MELLITUS WITH DIABETIC AUTONOMIC (POLY)NEUROPATHY|TYPE 1 DIABETES W DIABETIC AUTONOMIC (POLY)NEUROPATHY
C2874046|T047|E10.42|ICD10CM|TYPE 1 DIABETES MELLITUS WITH DIABETIC POLYNEUROPATHY|TYPE 1 DIABETES MELLITUS WITH DIABETIC NEURALGIA
C0837007|T047|E10.41|ICD10AM|TYPE 1 DIABETES MELLITUS WITH DIABETIC MONONEUROPATHY|TYPE 1 DIABETES MELLITUS WITH DIABETIC MONONEUROPATHY
C2874045|T047|E10.40|ICD10CM|TYPE 1 DIABETES MELLITUS WITH DIABETIC NEUROPATHY, UNSPECIFIED|TYPE 1 DIABETES MELLITUS WITH DIABETIC NEUROPATHY, UNSP
C2854087|T191|C91.00|ICD10CM|ACUTE LYMPHOBLASTIC LEUKEMIA NOT HAVING ACHIEVED REMISSION|ACUTE LYMPHOBLASTIC LEUKEMIA NOT HAVING ACHIEVED REMISSION
C0153876|T191||ICD10AM|ACUTE LYMPHOBLASTIC LEUKEMIA, IN REMISSION
C2854088|T191|C91.02|ICD10CM|ACUTE LYMPHOBLASTIC LEUKEMIA, IN RELAPSE|ACUTE LYMPHOBLASTIC LEUKEMIA, IN RELAPSE
C2874049|T047|E10.44|ICD10CM|TYPE 1 DIABETES MELLITUS WITH DIABETIC AMYOTROPHY|TYPE 1 DIABETES MELLITUS WITH DIABETIC AMYOTROPHY
C2890767|T037|T84.390A|ICD10CM|OTHER MECHANICAL COMPLICATION OF ELECTRONIC BONE STIMULATOR, INITIAL ENCOUNTER|MECH COMPL OF ELECTRONIC BONE STIMULATOR, INITIAL ENCOUNTER
C3263986|T047|G40.824|ICD10CM|EPILEPTIC SPASMS, INTRACTABLE, WITHOUT STATUS EPILEPTICUS|EPILEPTIC SPASMS, INTRACTABLE, WITHOUT STATUS EPILEPTICUS
C3263983|T047|G40.821|ICD10CM|EPILEPTIC SPASMS, NOT INTRACTABLE, WITH STATUS EPILEPTICUS|EPILEPTIC SPASMS, NOT INTRACTABLE, WITH STATUS EPILEPTICUS
C3263985|T047|G40.823|ICD10CM|EPILEPTIC SPASMS, INTRACTABLE, WITH STATUS EPILEPTICUS|EPILEPTIC SPASMS, INTRACTABLE, WITH STATUS EPILEPTICUS
C3263984|T047|G40.822|ICD10CM|EPILEPTIC SPASMS, NOT INTRACTABLE, WITHOUT STATUS EPILEPTICUS|EPILEPTIC SPASMS, NOT INTRACTABLE, W/O STATUS EPILEPTICUS
C4269550|T037|S02.670S|ICD10CM|FRACTURE OF ALVEOLUS OF MANDIBLE, UNSPECIFIED SIDE, SEQUELA|FRACTURE OF ALVEOLUS OF MANDIBLE, UNSPECIFIED SIDE, SEQUELA
C4269578|T037|S02.81XS|ICD10CM|FRACTURE OF OTHER SPECIFIED SKULL AND FACIAL BONES, RIGHT SIDE, SEQUELA|FRACTURE OF OTH SKULL AND FACIAL BONES, RIGHT SIDE, SEQUELA
C2835831|T037|S24.144D|ICD10CM|BROWN-SEQUARD SYNDROME AT T11-T12 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|BROWN-SEQUARD SYNDROME AT T11-T12, SUBS
C2833925|T037|S14.122S|ICD10CM|CENTRAL CORD SYNDROME AT C2 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|CENTRAL CORD SYNDROME AT C2, SEQUELA
C2835830|T037|S24.144A|ICD10CM|BROWN-SEQUARD SYNDROME AT T11-T12 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|BROWN-SEQUARD SYNDROME AT T11-T12, INIT
C2901847|T047|M86.329|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, UNSPECIFIED HUMERUS|CHRONIC MULTIFOCAL OSTEOMYELITIS, UNSPECIFIED HUMERUS
C4269574|T037|S02.81XB|ICD10CM|FRACTURE OF OTHER SPECIFIED SKULL AND FACIAL BONES, RIGHT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF OTH SKULL AND FACIAL BONES, RIGHT SIDE, 7THB
C4269573|T037|S02.81XA|ICD10CM|FRACTURE OF OTHER SPECIFIED SKULL AND FACIAL BONES, RIGHT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF OTH SKULL AND FACIAL BONES, RIGHT SIDE, INIT
C2901846|T047|M86.322|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, LEFT HUMERUS|CHRONIC MULTIFOCAL OSTEOMYELITIS, LEFT HUMERUS
C2833923|T037|S14.122A|ICD10CM|CENTRAL CORD SYNDROME AT C2 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|CENTRAL CORD SYNDROME AT C2, INIT
C2859215|T037|S73.032A|ICD10CM|OTHER ANTERIOR SUBLUXATION OF LEFT HIP, INITIAL ENCOUNTER|OTHER ANTERIOR SUBLUXATION OF LEFT HIP, INITIAL ENCOUNTER
C2901845|T047|M86.321|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, RIGHT HUMERUS|CHRONIC MULTIFOCAL OSTEOMYELITIS, RIGHT HUMERUS
C2833924|T037|S14.122D|ICD10CM|CENTRAL CORD SYNDROME AT C2 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|CENTRAL CORD SYNDROME AT C2, SUBS
C2835832|T037|S24.144S|ICD10CM|BROWN-SEQUARD SYNDROME AT T11-T12 LEVEL OF THORACIC SPINAL CORD, SEQUELA|BROWN-SEQUARD SYNDROME AT T11-T12, SEQUELA
C2855931|T037|S68.126S|ICD10CM|PARTIAL TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF RIGHT LITTLE FINGER, SEQUELA|PARTIAL TRAUMATIC MCP AMPUTATION OF R LITTLE FINGER, SEQUELA
C2882620|T047|I69.839|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING UNSPECIFIED SIDE|MONOPLG UPR LMB FOL OTH CEREBVASC DISEASE AFF UNSP SIDE
C2831503|T037|S02.413S|ICD10CM|LEFORT III FRACTURE, SEQUELA|LEFORT III FRACTURE, SEQUELA
C0338807|T048|F20.89|ICD10CM|OTHER SCHIZOPHRENIA|CENESTHOPATHIC SCHIZOPHRENIA
C2882616|T047|I69.831|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING RIGHT DOMINANT SIDE|MONOPLG UPR LMB FOL OTH CEREBVASC DISEASE AFF RIGHT DOM SIDE
C2882618|T047|I69.833|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING RIGHT NON-DOMINANT SIDE|MONOPLG UPR LMB FOL OTH CEREBVASC DIS AFF RIGHT NONDOM SIDE
C2882617|T047|I69.832|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING LEFT DOMINANT SIDE|MONOPLG UPR LMB FOL OTH CEREBVASC DISEASE AFF LEFT DOM SIDE
C0865304|T048||ICD10CM|SCHIZOPHRENIFORM DISORDER
C2882619|T047|I69.834|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING LEFT NON-DOMINANT SIDE|MONOPLG UPR LMB FOL OTH CEREBVASC DIS AFF LEFT NONDOM SIDE
C2831499|T037|S02.413B|ICD10CM|LEFORT III FRACTURE, INITIAL ENCOUNTER FOR OPEN FRACTURE|LEFORT III FRACTURE, INITIAL ENCOUNTER FOR OPEN FRACTURE
C2831498|T037|S02.413A|ICD10CM|LEFORT III FRACTURE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|LEFORT III FRACTURE, INITIAL ENCOUNTER FOR CLOSED FRACTURE
C2837905|T037|S32.409B|ICD10CM|UNSPECIFIED FRACTURE OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF UNSP ACETABULUM, INIT FOR OPN FX
C4270507|T046|T85.192A|ICD10CM|OTHER MECHANICAL COMPLICATION OF IMPLANTED ELECTRONIC NEUROSTIMULATOR OF SPINAL CORD ELECTRODE (LEAD), INITIAL ENCOUNTER|MECH COMPL OF IMPLNT ELEC NSTIM OF SPINAL CORD LEAD, INIT
C2857034|T037|S72.066B|ICD10CM|NONDISPLACED ARTICULAR FRACTURE OF HEAD OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP ARTIC FX HEAD OF UNSP FEMR, INIT FOR OPN FX TYPE I/2
C2890044|T037|T82.523A|ICD10CM|DISPLACEMENT OF BALLOON (COUNTERPULSATION) DEVICE, INITIAL ENCOUNTER|DISPLACEMENT OF BALLOON (COUNTERPULSATION) DEVICE, INIT
C0393517|T047|G32.81|ICD10CM|CEREBELLAR ATAXIA IN DISEASES CLASSIFIED ELSEWHERE|CEREBELLAR ATAXIA IN DISEASES CLASSIFIED ELSEWHERE
C2886765|T037|T79.A22A|ICD10CM|TRAUMATIC COMPARTMENT SYNDROME OF LEFT LOWER EXTREMITY, INITIAL ENCOUNTER|TRAUMATIC COMPARTMENT SYNDROME OF LEFT LOWER EXTREMITY, INIT
C2889233|T047|M05.411|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT SHOULDER|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF RIGHT SHOULDER
C4237245|T048|F11.94|ICD10CM|OPIOID USE, UNSPECIFIED WITH OPIOID-INDUCED MOOD DISORDER|OPIOID INDUCED DEPRESSIVE DISORDER, WITHOUT USE DISORDER
C2889234|T047|M05.412|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT SHOULDER|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF LEFT SHOULDER
C2874459|T048|F11.93|ICD10CM|OPIOID USE, UNSPECIFIED WITH WITHDRAWAL|OPIOID USE, UNSPECIFIED WITH WITHDRAWAL
C2889235|T047|M05.419|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF UNSP SHOULDER
C2874469|T048|F11.99|ICD10CM|OPIOID USE, UNSPECIFIED WITH UNSPECIFIED OPIOID-INDUCED DISORDER|OPIOID USE, UNSP WITH UNSPECIFIED OPIOID-INDUCED DISORDER
C2879364|T037|T45.92XS|ICD10CM|POISONING BY UNSPECIFIED PRIMARILY SYSTEMIC AND HEMATOLOGICAL AGENT, INTENTIONAL SELF-HARM, SEQUELA|POISN BY UNSP PRIM SYS AND HEMATOLOG AGENT, SLF-HRM, SEQUELA
C2901998|T046|M87.136|ICD10CM|OSTEONECROSIS DUE TO DRUGS OF UNSPECIFIED ULNA|OSTEONECROSIS DUE TO DRUGS OF UNSPECIFIED ULNA
C0268274|T047|E75.00|ICD10CM|GM2 GANGLIOSIDOSIS, UNSPECIFIED|GM2 GANGLIOSIDOSIS, UNSPECIFIED
C0036161|T047||ICD10CM|SANDHOFF DISEASE
C0039373|T047||ICD10CM|TAY-SACHS DISEASE
C1527407|T047||ICD10CM|PULMONARY EOSINOPHILIA, NOT ELSEWHERE CLASSIFIED
C2874271|T047|E75.09|ICD10CM|OTHER GM2 GANGLIOSIDOSIS|OTHER GM2 GANGLIOSIDOSIS
C2901488|T046|M84.652A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, LEFT FEMUR, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, LEFT FEMUR, INIT
C2856551|T037|S72.012A|ICD10CM|UNSPECIFIED INTRACAPSULAR FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP INTRACAPSULAR FRACTURE OF LEFT FEMUR, INIT FOR CLOS FX
C2856552|T037|S72.012B|ICD10CM|UNSPECIFIED INTRACAPSULAR FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP INTRACAP FX LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C2876693|T037|T36.6X2A|ICD10CM|POISONING BY RIFAMPICINS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY RIFAMPICINS, INTENTIONAL SELF-HARM, INIT ENCNTR
C2884929|T037|T59.6X2A|ICD10CM|TOXIC EFFECT OF HYDROGEN SULFIDE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF HYDROGEN SULFIDE, SELF-HARM, INIT
C2880089|T047|A01.04|ICD10CM|TYPHOID ARTHRITIS|TYPHOID ARTHRITIS
C2856553|T037|S72.012C|ICD10CM|UNSPECIFIED INTRACAPSULAR FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP INTRACAP FX LEFT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2977000|T046|I82.4Z9|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF UNSPECIFIED DISTAL LOWER EXTREMITY|ACUTE EMBLSM AND THOMBOS UNSP DEEP VN UNSP DISTAL LOW EXTRM
C2858374|T037|S72.413C|ICD10CM|DISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL UNSP CONDYLE FX LOW END UNSP FEMR, 7THC
C2833621|T037|S12.650A|ICD10CM|OTHER TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH TRAUM DISPL SPONDYLOLYSIS OF SEVENTH CERVCAL VERT, INIT
C2858373|T037|S72.413B|ICD10CM|DISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL UNSP CONDYLE FX LOW END UNSP FEMR, 7THB
C2976997|T046|I82.4Z1|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF RIGHT DISTAL LOWER EXTREMITY|AC EMBLSM AND THOMBOS UNSP DEEP VEINS OF R DIST LOW EXTRM
C2976999|T046|I82.4Z3|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF DISTAL LOWER EXTREMITY, BILATERAL|AC EMBLSM AND THOMBOS UNSP DEEP VEINS OF DIST LOW EXTRM, BI
C2976998|T046|I82.4Z2|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF LEFT DISTAL LOWER EXTREMITY|AC EMBLSM AND THOMBOS UNSP DEEP VEINS OF LEFT DIST LOW EXTRM
C2858372|T037|S72.413A|ICD10CM|DISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED UNSP CONDYLE FX LOWER END OF UNSP FEMUR, INIT
C2890887|T037|T84.63XA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL FIXATION DEVICE OF SPINE, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INT FIX OF SPINE, INIT
C2838515|T037|S32.9XXA|ICD10CM|FRACTURE OF UNSPECIFIED PARTS OF LUMBOSACRAL SPINE AND PELVIS, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF UNSP PARTS OF LUMBOSACRAL SPINE AND PELVIS, INIT
C2838516|T037|S32.9XXB|ICD10CM|FRACTURE OF UNSPECIFIED PARTS OF LUMBOSACRAL SPINE AND PELVIS, INITIAL ENCOUNTER FOR OPEN FRACTURE|FX UNSP PARTS OF LUMBOSACRAL SPINE & PELVIS, INIT FOR OPN FX
C2830415|T033|R40.2324|ICD10CM|COMA SCALE, BEST MOTOR RESPONSE, EXTENSION, 24 HOURS OR MORE AFTER HOSPITAL ADMISSION|COMA SCALE, BEST MOTOR RESPONSE, EXTENSION, 24+HRS
C2876643|T037|T36.4X2A|ICD10CM|POISONING BY TETRACYCLINES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY TETRACYCLINES, INTENTIONAL SELF-HARM, INIT
C2830413|T033|R40.2322|ICD10CM|COMA SCALE, BEST MOTOR RESPONSE, EXTENSION, AT ARRIVAL TO EMERGENCY DEPARTMENT|COMA SCALE, BEST MOTOR RESPONSE, EXTENSION, EMR
C2830414|T033|R40.2323|ICD10CM|COMA SCALE, BEST MOTOR RESPONSE, EXTENSION, AT HOSPITAL ADMISSION|COMA SCALE, BEST MOTOR RESPONSE, EXTENSION, ADMIT
C2830411|T033|R40.2320|ICD10CM|COMA SCALE, BEST MOTOR RESPONSE, EXTENSION, UNSPECIFIED TIME|COMA SCALE, BEST MOTOR RESPONSE, EXTENSION, UNSPECIFIED TIME
C2830412|T033|R40.2321|ICD10CM|COMA SCALE, BEST MOTOR RESPONSE, EXTENSION, IN THE FIELD [EMT OR AMBULANCE]|COMA SCALE, BEST MOTOR RESPONSE, EXTENSION, IN THE FIELD
C4268026|T047|E10.3399|ICD10CM|TYPE 1 DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|TYPE 1 DIAB WITH MOD NONP RTNOP WITHOUT MACULAR EDEMA, UNSP
C4268023|T047|E10.3391|ICD10CM|TYPE 1 DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|TYPE 1 DIAB WITH MOD NONP RTNOP WITHOUT MACULAR EDEMA, R EYE
C4268024|T047|E10.3392|ICD10CM|TYPE 1 DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|TYPE 1 DIAB WITH MOD NONP RTNOP WITHOUT MACULAR EDEMA, L EYE
C4268025|T047|E10.3393|ICD10CM|TYPE 1 DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|TYPE 1 DIAB WITH MOD NONP RTNOP WITHOUT MACULAR EDEMA, BI
C2902735|T037|M96.65|ICD10CM|FRACTURE OF PELVIS FOLLOWING INSERTION OF ORTHOPEDIC IMPLANT, JOINT PROSTHESIS, OR BONE PLATE|FX PELVIS FOLLOWING INSRT ORTHO IMPLNT/PROSTH/BONE PLT
C2902744|T037|M96.69|ICD10CM|FRACTURE OF OTHER BONE FOLLOWING INSERTION OF ORTHOPEDIC IMPLANT, JOINT PROSTHESIS, OR BONE PLATE|FX BONE FOLLOWING INSRT ORTHO IMPLNT/PROSTH/BONE PLT
C0477405|T047|G72.89|ICD10CM|OTHER SPECIFIED MYOPATHIES|OTHER SPECIFIED MYOPATHIES
C2884947|T037|T59.7X2S|ICD10CM|TOXIC EFFECT OF CARBON DIOXIDE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CARBON DIOXIDE, SELF-HARM, SEQUELA
C1135346|T047|G72.81|ICD10CM|CRITICAL ILLNESS MYOPATHY|INTENSIVE CARE (ICU) MYOPATHY
C2855881|T037|S68.114S|ICD10CM|COMPLETE TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF RIGHT RING FINGER, SEQUELA|COMPLETE TRAUMATIC MCP AMPUTATION OF R RNG FNGR, SEQUELA
C1456240|T047|G47.419|ICD10CM|NARCOLEPSY WITHOUT CATAPLEXY|NARCOLEPSY WITHOUT CATAPLEXY
C2902079|T046|M87.279|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED TOE(S)|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED TOE(S)
C2902078|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, LEFT TOE(S)
C2902077|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, RIGHT TOE(S)
C2902076|T046|M87.276|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED FOOT|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED FOOT
C2902075|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, LEFT FOOT
C2902074|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, RIGHT FOOT
C0751362|T047||ICD10CM|NARCOLEPSY WITH CATAPLEXY
C2902072|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, LEFT ANKLE
C2902071|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, RIGHT ANKLE
C4270326|T046|T83.518A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO OTHER URINARY CATHETER, INITIAL ENCOUNTER|I/I REACT D/T OTHER URINARY CATHETER, INITIAL ENCOUNTER
C2882086|T047|I13.2|ICD10CM|HYPERTENSIVE HEART AND CHRONIC KIDNEY DISEASE WITH HEART FAILURE AND WITH STAGE 5 CHRONIC KIDNEY DISEASE, OR END STAGE RENAL DISEASE|HYP HRT & CHR KDNY DIS W HRT FAIL AND W STG 5 CHR KDNY/ESRD
C2882081|T047|I13.0|ICD10CM|HYPERTENSIVE HEART AND CHRONIC KIDNEY DISEASE WITH HEART FAILURE AND STAGE 1 THROUGH STAGE 4 CHRONIC KIDNEY DISEASE, OR UNSPECIFIED CHRONIC KIDNEY DISEASE|HYP HRT & CHR KDNY DIS W HRT FAIL AND STG 1-4/UNSP CHR KDNY
C2890813|T037|T84.53XA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL RIGHT KNEE PROSTHESIS, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INTERNAL R KNEE PROSTH, INIT
C2845916|T191|C69.52|ICD10CM|MALIGNANT NEOPLASM OF LEFT LACRIMAL GLAND AND DUCT|MALIGNANT NEOPLASM OF LEFT LACRIMAL GLAND AND DUCT
C2905681|T037|X73.1XXS|ICD10CM|INTENTIONAL SELF-HARM BY HUNTING RIFLE DISCHARGE, SEQUELA|INTENTIONAL SELF-HARM BY HUNTING RIFLE DISCHARGE, SEQUELA
C2845914|T191|C69.50|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED LACRIMAL GLAND AND DUCT|MALIGNANT NEOPLASM OF UNSPECIFIED LACRIMAL GLAND AND DUCT
C2845915|T191|C69.51|ICD10CM|MALIGNANT NEOPLASM OF RIGHT LACRIMAL GLAND AND DUCT|MALIGNANT NEOPLASM OF RIGHT LACRIMAL GLAND AND DUCT
C2879078|T037|T45.2X2S|ICD10CM|POISONING BY VITAMINS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY VITAMINS, INTENTIONAL SELF-HARM, SEQUELA
C2889430|T047|M06.259|ICD10CM|RHEUMATOID BURSITIS, UNSPECIFIED HIP|RHEUMATOID BURSITIS, UNSPECIFIED HIP
C2882379|T047|I63.39|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF OTHER CEREBRAL ARTERY|CEREBRAL INFARCTION DUE TO THROMBOSIS OF OTH CEREBRAL ARTERY
C2889429|T047|M06.252|ICD10CM|RHEUMATOID BURSITIS, LEFT HIP|RHEUMATOID BURSITIS, LEFT HIP
C2889428|T047|M06.251|ICD10CM|RHEUMATOID BURSITIS, RIGHT HIP|RHEUMATOID BURSITIS, RIGHT HIP
C2879103|T037|T45.3X2S|ICD10CM|POISONING BY ENZYMES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ENZYMES, INTENTIONAL SELF-HARM, SEQUELA
C2888029|T046|K94.19|ICD10CM|OTHER COMPLICATIONS OF ENTEROSTOMY|OTHER COMPLICATIONS OF ENTEROSTOMY
C1443975|T047|K94.12|ICD10CM|ENTEROSTOMY INFECTION|ENTEROSTOMY INFECTION
C2118344|T046|K94.13|ICD10CM|ENTEROSTOMY MALFUNCTION|MECHANICAL COMPLICATION OF ENTEROSTOMY
C2888027|T046|K94.10|ICD10CM|ENTEROSTOMY COMPLICATION, UNSPECIFIED|ENTEROSTOMY COMPLICATION, UNSPECIFIED
C2888028|T046|K94.11|ICD10CM|ENTEROSTOMY HEMORRHAGE|ENTEROSTOMY HEMORRHAGE
C2879101|T037|T45.3X2A|ICD10CM|POISONING BY ENZYMES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ENZYMES, INTENTIONAL SELF-HARM, INIT ENCNTR
C2889482|T047|M06.851|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, RIGHT HIP|OTHER SPECIFIED RHEUMATOID ARTHRITIS, RIGHT HIP
C2889483|T047|M06.852|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, LEFT HIP|OTHER SPECIFIED RHEUMATOID ARTHRITIS, LEFT HIP
C2889448|T046|M06.331|ICD10CM|RHEUMATOID NODULE, RIGHT WRIST|RHEUMATOID NODULE, RIGHT WRIST
C2889449|T046|M06.332|ICD10CM|RHEUMATOID NODULE, LEFT WRIST|RHEUMATOID NODULE, LEFT WRIST
C2889450|T046|M06.339|ICD10CM|RHEUMATOID NODULE, UNSPECIFIED WRIST|RHEUMATOID NODULE, UNSPECIFIED WRIST
C2890433|T037|T84.021A|ICD10CM|DISLOCATION OF INTERNAL LEFT HIP PROSTHESIS, INITIAL ENCOUNTER|DISLOCATION OF INTERNAL LEFT HIP PROSTHESIS, INIT ENCNTR
C2977877|T037|S32.599B|ICD10CM|OTHER SPECIFIED FRACTURE OF UNSPECIFIED PUBIS, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF UNSP PUBIS, INIT ENCNTR FOR OPEN FRACTURE
C2838423|T037|S32.609B|ICD10CM|UNSPECIFIED FRACTURE OF UNSPECIFIED ISCHIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF UNSP ISCHIUM, INIT ENCNTR FOR OPEN FRACTURE
C2837567|T037|S32.032A|ICD10CM|UNSTABLE BURST FRACTURE OF THIRD LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSTABLE BURST FRACTURE OF THIRD LUMBAR VERTEBRA, INIT
C2874848|T048|F19.951|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH PSYCHOACTIVE SUBSTANCE-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|OTH PSYCHOACTV SUB USE, UNSP W PSYCH DISORDER W HALLUCIN
C0349354|T191|C43.8|DMDICD10|MALIGNANT MELANOMA OF OVERLAPPING SITES OF SKIN|BOESARTIGES MELANOM DER HAUT, MEHRERE TEILBEREICHE UEBERLAPPEND
C2977901|T191|C43.9|ICD10CM|MALIGNANT MELANOMA OF SKIN, UNSPECIFIED|MALIGNANT MELANOMA OF UNSPECIFIED SITE OF SKIN
C2901010|T046|M84.454A|ICD10CM|PATHOLOGICAL FRACTURE, PELVIS, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, PELVIS, INIT ENCNTR FOR FRACTURE
C0153529|T191|C43.0|DMDICD10|MALIGNANT MELANOMA OF LIP|BOESARTIGES MELANOM DER LIPPE
C0346782|T191|C43.4|DMDICD10|MALIGNANT MELANOMA OF SCALP AND NECK|BOESARTIGES MELANOM DER BEHAARTEN KOPFHAUT UND DES HALSES
C2869774|T037|S98.022S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT FOOT AT ANKLE LEVEL, SEQUELA|PARTIAL TRAUMATIC AMP OF LEFT FOOT AT ANKLE LEVEL, SEQUELA
C2889943|T037|T82.332A|ICD10CM|LEAKAGE OF FEMORAL ARTERIAL GRAFT (BYPASS), INITIAL ENCOUNTER|LEAKAGE OF FEMORAL ARTERIAL GRAFT (BYPASS), INIT ENCNTR
C0037899|T047|E75.3|DMDICD10|SPHINGOLIPIDOSIS, UNSPECIFIED|SPHINGOLIPIDOSE, NICHT NAEHER BEZEICHNET
C0342342|T047|E20.0|DMDICD10|IDIOPATHIC HYPOPARATHYROIDISM|IDIOPATHISCHER HYPOPARATHYREOIDISMUS
C0023794|T047|E75.6|DMDICD10|LIPID STORAGE DISORDER, UNSPECIFIED|STOERUNG DER LIPIDSPEICHERUNG, NICHT NAEHER BEZEICHNET
C2874275|T047|E75.5|ICD10CM|OTHER LIPID STORAGE DISORDERS|CEREBROTENDINOUS CHOLESTEROSIS [VAN BOGAERT-SCHERER-EPSTEIN]
C0751383|T047||ICD10CM|NEURONAL CEROID LIPOFUSCINOSIS
C0242037|T047||ICD10CM|HYPOPARATHYROIDISM, UNSPECIFIED
C0348454|T047|E20.8|DMDICD10|OTHER HYPOPARATHYROIDISM|SONSTIGER HYPOPARATHYREOIDISMUS
C2832305|T037|S06.360A|ICD10CM|TRAUMATIC HEMORRHAGE OF CEREBRUM, UNSPECIFIED, WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|TRAUM HEMOR CEREB, W/O LOSS OF CONSCIOUSNESS, INIT
C2885156|T037|T61.772A|ICD10CM|OTHER FISH POISONING, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|OTHER FISH POISONING, INTENTIONAL SELF-HARM, INIT ENCNTR
C2888431|T047|L89.311|ICD10CM|PRESSURE ULCER OF RIGHT BUTTOCK, STAGE 1|PRESSURE ULCER OF RIGHT BUTTOCK, STAGE 1
C2888428|T047||ICD10CM|PRESSURE ULCER OF RIGHT BUTTOCK, UNSTAGEABLE
C2888437|T047|L89.313|ICD10CM|PRESSURE ULCER OF RIGHT BUTTOCK, STAGE 3|PRESSURE ULCER OF RIGHT BUTTOCK, STAGE 3
C2888434|T047|L89.312|ICD10CM|PRESSURE ULCER OF RIGHT BUTTOCK, STAGE 2|PRESSURE ULCER OF RIGHT BUTTOCK, STAGE 2
C2888440|T047|L89.314|ICD10CM|PRESSURE ULCER OF RIGHT BUTTOCK, STAGE 4|PRESSURE ULCER OF RIGHT BUTTOCK, STAGE 4
C4270481|T046|T85.121A|ICD10CM|DISPLACEMENT OF IMPLANTED ELECTRONIC NEUROSTIMULATOR OF PERIPHERAL NERVE ELECTRODE (LEAD), INITIAL ENCOUNTER|DISPLACEMENT OF IMPLNT ELEC NSTIM OF PRPH NRV LEAD, INIT
C2888443|T047|L89.319|ICD10CM|PRESSURE ULCER OF RIGHT BUTTOCK, UNSPECIFIED STAGE|PRESSURE ULCER OF RIGHT BUTTOCK, UNSPECIFIED STAGE
C2832307|T037|S06.360S|ICD10CM|TRAUMATIC HEMORRHAGE OF CEREBRUM, UNSPECIFIED, WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|TRAUM HEMOR CEREB, W/O LOSS OF CONSCIOUSNESS, SEQUELA
C2885158|T037|T61.772S|ICD10CM|OTHER FISH POISONING, INTENTIONAL SELF-HARM, SEQUELA|OTHER FISH POISONING, INTENTIONAL SELF-HARM, SEQUELA
C2876151|T037|T31.63|ICD10CM|BURNS INVOLVING 60-69% OF BODY SURFACE WITH 30-39% THIRD DEGREE BURNS|BURNS OF 60-69% OF BODY SURFACE W 30-39% THIRD DEGREE BURNS
C4269377|T037|S02.40AA|ICD10CM|MALAR FRACTURE, RIGHT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|MALAR FRACTURE, RIGHT SIDE, INIT
C2882579|T047|I69.339|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING CEREBRAL INFARCTION AFFECTING UNSPECIFIED SIDE|MONOPLG UPR LMB FOLLOWING CEREBRAL INFRC AFFECTING UNSP SIDE
C2882578|T047|I69.334|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING CEREBRAL INFARCTION AFFECTING LEFT NON-DOMINANT SIDE|MONOPLG UPR LMB FOL CEREBRAL INFRC AFF LEFT NONDOM SIDE
C2832364|T037|S06.374S|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF CEREBELLUM WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|CONTUS/LAC/HEM CRBLM W LOC OF 6 HOURS TO 24 HOURS, SEQUELA
C2882576|T047|I69.332|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING CEREBRAL INFARCTION AFFECTING LEFT DOMINANT SIDE|MONOPLG UPR LMB FOL CEREBRAL INFRC AFF LEFT DOMINANT SIDE
C2882577|T047|I69.333|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING CEREBRAL INFARCTION AFFECTING RIGHT NON-DOMINANT SIDE|MONOPLG UPR LMB FOL CEREBRAL INFRC AFF RIGHT NONDOM SIDE
C2882575|T047|I69.331|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING CEREBRAL INFARCTION AFFECTING RIGHT DOMINANT SIDE|MONOPLG UPR LMB FOL CEREBRAL INFRC AFF RIGHT DOMINANT SIDE
C2893390|T047|A54.43|ICD10CM|GONOCOCCAL OSTEOMYELITIS|GONOCOCCAL OSTEOMYELITIS
C0153216|T047|A54.42|ICD10CM|GONOCOCCAL ARTHRITIS|GONOCOCCAL ARTHRITIS
C2893389|T047|A54.41|ICD10CM|GONOCOCCAL SPONDYLOPATHY|GONOCOCCAL SPONDYLOPATHY
C0494057|T047|A54.40|ICD10CM|GONOCOCCAL INFECTION OF MUSCULOSKELETAL SYSTEM, UNSPECIFIED|GONOCOCCAL INFECTION OF MUSCULOSKELETAL SYSTEM, UNSPECIFIED
C2832362|T037|S06.374A|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF CEREBELLUM WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|CONTUS/LAC/HEM CRBLM W LOC OF 6 HOURS TO 24 HOURS, INIT
C4269305|T037|S02.11DS|ICD10CM|TYPE II OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, SEQUELA|TYPE II OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, SEQUELA
C1719298|T047|B00.82|ICD10CM|HERPES SIMPLEX MYELITIS|HERPES SIMPLEX MYELITIS
C2893392|T047|A54.49|ICD10CM|GONOCOCCAL INFECTION OF OTHER MUSCULOSKELETAL TISSUE|GONOCOCCAL INFECTION OF OTHER MUSCULOSKELETAL TISSUE
C2876150|T037|T31.62|ICD10CM|BURNS INVOLVING 60-69% OF BODY SURFACE WITH 20-29% THIRD DEGREE BURNS|BURNS OF 60-69% OF BODY SURFACE W 20-29% THIRD DEGREE BURNS
C2900518|T046|M80.859A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, UNSP FEMUR, INIT
C2889008|T047|M02.149|ICD10CM|POSTDYSENTERIC ARTHROPATHY, UNSPECIFIED HAND|POSTDYSENTERIC ARTHROPATHY, UNSPECIFIED HAND
C2885577|T037|T63.332S|ICD10CM|TOXIC EFFECT OF VENOM OF BROWN RECLUSE SPIDER, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF BROWN RECLUSE SPIDER, SLF-HRM, SQLA
C4268611|T047|K55.011|ICD10CM|FOCAL (SEGMENTAL) ACUTE (REVERSIBLE) ISCHEMIA OF SMALL INTESTINE|FOCAL (SEGMENTAL) ACUTE ISCHEMIA OF SMALL INTESTINE
C2889007|T047|M02.142|ICD10CM|POSTDYSENTERIC ARTHROPATHY, LEFT HAND|POSTDYSENTERIC ARTHROPATHY, LEFT HAND
C2889006|T047|M02.141|ICD10CM|POSTDYSENTERIC ARTHROPATHY, RIGHT HAND|POSTDYSENTERIC ARTHROPATHY, RIGHT HAND
C2837981|T191|C40.82|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF BONE AND ARTICULAR CARTILAGE OF LEFT LIMB|MALIG NEOPLM OF OVRLP SITES OF BONE/ARTIC CARTL OF LEFT LIMB
C2837979|T191|C40.80|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF BONE AND ARTICULAR CARTILAGE OF UNSPECIFIED LIMB|MALIG NEOPLM OF OVRLP SITES OF BONE/ARTIC CARTL OF UNSP LIMB
C2837980|T191|C40.81|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF BONE AND ARTICULAR CARTILAGE OF RIGHT LIMB|MALIG NEOPLM OF OVRLP SITES OF BONE/ARTIC CARTL OF R LIMB
C2890618|T037|T84.120A|ICD10CM|DISPLACEMENT OF INTERNAL FIXATION DEVICE OF RIGHT HUMERUS, INITIAL ENCOUNTER|DISPLACEMENT OF INT FIX OF RIGHT HUMERUS, INIT
C2885575|T037|T63.332A|ICD10CM|TOXIC EFFECT OF VENOM OF BROWN RECLUSE SPIDER, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF BROWN RECLUSE SPIDER, SLF-HRM, INIT
C2902439|T047|M90.549|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, UNSPECIFIED HAND|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, UNSP HAND
C2882509|T047|I69.159|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING UNSPECIFIED SIDE|HEMIPLGA FOLLOWING NTRM INTCRBL HEMOR AFFECTING UNSP SIDE
C2882506|T047|I69.152|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING LEFT DOMINANT SIDE|HEMIPLGA FOLLOWING NTRM INTCRBL HEMOR AFF LEFT DOMINANT SIDE
C2882507|T047|I69.153|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING RIGHT NON-DOMINANT SIDE|HEMIPLGA FOLLOWING NTRM INTCRBL HEMOR AFF RIGHT NONDOM SIDE
C2882505|T047|I69.151|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING RIGHT DOMINANT SIDE|HEMIPLGA FOL NTRM INTCRBL HEMOR AFF RIGHT DOMINANT SIDE
C2873865|T047|E05.01|ICD10CM|THYROTOXICOSIS WITH DIFFUSE GOITER WITH THYROTOXIC CRISIS OR STORM|THYROTOXICOSIS W DIFFUSE GOITER W THYROTOXIC CRISIS OR STORM
C2873864|T047|E05.00|ICD10CM|THYROTOXICOSIS WITH DIFFUSE GOITER WITHOUT THYROTOXIC CRISIS OR STORM|THYROTOXICOSIS W DIFFUSE GOITER W/O THYROTOXIC CRISIS
C2882508|T047|I69.154|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING LEFT NON-DOMINANT SIDE|HEMIPLGA FOLLOWING NTRM INTCRBL HEMOR AFF LEFT NONDOM SIDE
C2874721|T048|F16.99|ICD10CM|HALLUCINOGEN USE, UNSPECIFIED WITH UNSPECIFIED HALLUCINOGEN-INDUCED DISORDER|HALLUCINOGEN USE, UNSP W UNSP HALLUCINOGEN-INDUCED DISORDER
C2902954|T047|N17.2|ICD10CM|ACUTE KIDNEY FAILURE WITH MEDULLARY NECROSIS|RENAL MEDULLARY [PAPILLARY] NECROSIS
C2858216|T037|S72.366A|ICD10CM|NONDISPLACED SEGMENTAL FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED SEGMENTAL FRACTURE OF SHAFT OF UNSP FEMUR, INIT
C4268274|T048|F16.94|ICD10CM|HALLUCINOGEN USE, UNSPECIFIED WITH HALLUCINOGEN-INDUCED MOOD DISORDER|PHENCYCLIDINE INDUCED BIPOLAR OR RELATED DISORDER, WITHOUT USE DISORDER
C2838678|T037|S34.124A|ICD10CM|INCOMPLETE LESION OF L4 LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|INCOMPLETE LESION OF L4 LEVEL OF LUMBAR SPINAL CORD, INIT
C0348495|T047|E78.8|ICD10CM|OTHER LIPOPROTEIN METABOLISM DISORDERS|OTHER DISORDERS OF LIPOPROTEIN METABOLISM
C2887151|T047|I82.B19|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED SUBCLAVIAN VEIN|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED SUBCLAVIAN VEIN
C0311284|T047|E78.81|ICD10CM|LIPOID DERMATOARTHRITIS|LIPOID DERMATOARTHRITIS
C2887150|T047|I82.B13|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF SUBCLAVIAN VEIN, BILATERAL|ACUTE EMBOLISM AND THROMBOSIS OF SUBCLAVIAN VEIN, BILATERAL
C2833286|T037|S12.150A|ICD10CM|OTHER TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH TRAUM DISPL SPONDYLOLYSIS OF SECOND CERVCAL VERT, INIT
C2887148|T047|I82.B11|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF RIGHT SUBCLAVIAN VEIN|ACUTE EMBOLISM AND THROMBOSIS OF RIGHT SUBCLAVIAN VEIN
C2901890|T047|M86.511|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, RIGHT SHOULDER|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, RIGHT SHOULDER
C2857412|T037|S72.134B|ICD10CM|NONDISPLACED APOPHYSEAL FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP APOPHYSEAL FX RIGHT FEMUR, INIT FOR OPN FX TYPE I/2
C2857411|T037|S72.134A|ICD10CM|NONDISPLACED APOPHYSEAL FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED APOPHYSEAL FRACTURE OF RIGHT FEMUR, INIT
C2901891|T047|M86.512|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, LEFT SHOULDER|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, LEFT SHOULDER
C2901892|T047|M86.51|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED SHOULDER|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, SHOULDER
C2875158|T047|G43.411|ICD10CM|HEMIPLEGIC MIGRAINE, INTRACTABLE, WITH STATUS MIGRAINOSUS|HEMIPLEGIC MIGRAINE, INTRACTABLE, WITH STATUS MIGRAINOSUS
C4268255|T048|F15.24|ICD10CM|OTHER STIMULANT DEPENDENCE WITH STIMULANT-INDUCED MOOD DISORDER|AMPHETAMINE OR OTHER STIMULANT USE DISORDER, SEVERE, WITH AMPHETAMINE OR OTHER STIMULANT-INDUCED DEPRESSIVE DISORDER
C4236987|T048|F15.23|ICD10CM|OTHER STIMULANT DEPENDENCE WITH WITHDRAWAL|AMPHETAMINE OR OTHER STIMULANT WITHDRAWAL
C2838236|T037|S32.463A|ICD10CM|DISPLACED ASSOCIATED TRANSVERSE-POSTERIOR FRACTURE OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED ASSOCIATED TRANSV/POST FX UNSP ACETABULUM, INIT
C4509067|T048|F15.21|ICD10CM|OTHER STIMULANT DEPENDENCE, IN REMISSION|AMPHETAMINE TYPE SUBSTANCE USE DISORDER, SEVERE, IN SUSTAINED REMISSION
C4237318|T048|F15.20|ICD10CM|OTHER STIMULANT DEPENDENCE, UNCOMPLICATED|OTHER OR UNSPECIFIED STIMULANT USE DISORDER, SEVERE
C2875159|T047|G43.419|ICD10CM|HEMIPLEGIC MIGRAINE, INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|HEMIPLEGIC MIGRAINE, INTRACTABLE, WITHOUT STATUS MIGRAINOSUS
C4269515|T037|S02.641S|ICD10CM|FRACTURE OF RAMUS OF RIGHT MANDIBLE, SEQUELA|FRACTURE OF RAMUS OF RIGHT MANDIBLE, SEQUELA
C2884253|T037|T53.3X2A|ICD10CM|TOXIC EFFECT OF TETRACHLOROETHYLENE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF TETRACHLOROETHYLENE, SELF-HARM, INIT
C2874660|T048|F15.29|ICD10CM|OTHER STIMULANT DEPENDENCE WITH UNSPECIFIED STIMULANT-INDUCED DISORDER|OTH STIMULANT DEPENDENCE W UNSP STIMULANT-INDUCED DISORDER
C2890756|T037|T84.320A|ICD10CM|DISPLACEMENT OF ELECTRONIC BONE STIMULATOR, INITIAL ENCOUNTER|DISPLACEMENT OF ELECTRONIC BONE STIMULATOR, INIT ENCNTR
C2874029|T047|E10.311|ICD10CM|TYPE 1 DIABETES MELLITUS WITH UNSPECIFIED DIABETIC RETINOPATHY WITH MACULAR EDEMA|TYPE 1 DIABETES W UNSP DIABETIC RETINOPATHY W MACULAR EDEMA
C2856007|T037|S68.611S|ICD10CM|COMPLETE TRAUMATIC TRANSPHALANGEAL AMPUTATION OF LEFT INDEX FINGER, SEQUELA|COMPLETE TRAUMATIC TRNSPHAL AMP OF L IDX FNGR, SEQUELA
C2349570|T037||ICD10CM|ACUTE KIDNEY FAILURE, UNSPECIFIED
C2874030|T047|E10.319|ICD10CM|TYPE 1 DIABETES MELLITUS WITH UNSPECIFIED DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA|TYPE 1 DIABETES W UNSP DIABETIC RTNOP W/O MACULAR EDEMA
C2884255|T037|T53.3X2S|ICD10CM|TOXIC EFFECT OF TETRACHLOROETHYLENE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF TETRACHLOROETHYLENE, SELF-HARM, SEQUELA
C4087321|T048|F45.1|ICD10CM|UNDIFFERENTIATED SOMATOFORM DISORDER|SOMATIC SYMPTOM DISORDER
C1405656|T048||ICD10CM|SOMATIZATION DISORDER
C2838643|T037|S34.111S|ICD10CM|COMPLETE LESION OF L1 LEVEL OF LUMBAR SPINAL CORD, SEQUELA|COMPLETE LESION OF L1 LEVEL OF LUMBAR SPINAL CORD, SEQUELA
C0037650|T048|F45|DMDICD10|SOMATOFORM DISORDER, UNSPECIFIED|SOMATOFORME STOERUNGEN
C2874956|T048|F45.8|ICD10CM|OTHER SOMATOFORM DISORDERS|PSYCHOGENIC DYSPHAGIA, INCLUDING 'GLOBUS HYSTERICUS'
C0036391|T047|G71.13|ICD10CM|MYOTONIC CHONDRODYSTROPHY|SCHWARTZ-JAMPEL DISEASE
C2936781|T047|G71.12|ICD10CM|MYOTONIA CONGENITA|DOMINANT MYOTONIA CONGENITA [THOMSEN DISEASE]
C1404542|T046||ICD10CM|DRUG INDUCED MYOTONIA
C2833856|T037|S14.103S|ICD10CM|UNSPECIFIED INJURY AT C3 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|UNSP INJURY AT C3 LEVEL OF CERVICAL SPINAL CORD, SEQUELA
C2882329|T047|I63.00|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF UNSPECIFIED PRECEREBRAL ARTERY|CEREBRAL INFARCTION DUE TO THOMBOS UNSP PRECEREBRAL ARTERY
C2882334|T047|I63.02|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF BASILAR ARTERY|CEREBRAL INFARCTION DUE TO THROMBOSIS OF BASILAR ARTERY
C2882339|T047|I63.09|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF OTHER PRECEREBRAL ARTERY|CEREBRAL INFARCTION DUE TO THROMBOSIS OF PRECEREBRAL ARTERY
C2833855|T037|S14.103D|ICD10CM|UNSPECIFIED INJURY AT C3 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY AT C3 LEVEL OF CERVICAL SPINAL CORD, SUBS ENCNTR
C2833854|T037|S14.103A|ICD10CM|UNSPECIFIED INJURY AT C3 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY AT C3 LEVEL OF CERVICAL SPINAL CORD, INIT ENCNTR
C2876745|T037|T36.8X2S|ICD10CM|POISONING BY OTHER SYSTEMIC ANTIBIOTICS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH SYSTEMIC ANTIBIOTICS, SELF-HARM, SEQUELA
C3161096|T047||ICD10CM|RESPIRATORY CONDITIONS DUE TO SMOKE INHALATION
C0348822|T046|J70.4|DMDICD10|DRUG-INDUCED INTERSTITIAL LUNG DISORDERS, UNSPECIFIED|ARZNEIMITTELINDUZIERTE INTERSTITIELLE LUNGENKRANKHEIT, NICHT NAEHER BEZEICHNET
C0340126|T047|J70.1|ICD10CM|CHRONIC AND OTHER PULMONARY MANIFESTATIONS DUE TO RADIATION|FIBROSIS OF LUNG FOLLOWING RADIATION
C0206063|T037||ICD10CM|ACUTE PULMONARY MANIFESTATIONS DUE TO RADIATION
C0348824|T046|J70.3|DMDICD10|CHRONIC DRUG-INDUCED INTERSTITIAL LUNG DISORDERS|CHRONISCHE ARZNEIMITTELINDUZIERTE INTERSTITIELLE LUNGENKRANKHEITEN
C0348823|T046|J70.2|DMDICD10|ACUTE DRUG-INDUCED INTERSTITIAL LUNG DISORDERS|AKUTE ARZNEIMITTELINDUZIERTE INTERSTITIELLE LUNGENKRANKHEITEN
C0155905|T047|J70.9|DMDICD10|RESPIRATORY CONDITIONS DUE TO UNSPECIFIED EXTERNAL AGENT|KRANKHEITEN DER ATMUNGSORGANE DURCH NICHT NAEHER BEZEICHNETE EXOGENE SUBSTANZ
C0155904|T047|J70.8|DMDICD10|RESPIRATORY CONDITIONS DUE TO OTHER SPECIFIED EXTERNAL AGENTS|KRANKHEITEN DER ATMUNGSORGANE DURCH SONSTIGE NAEHER BEZEICHNETE EXOGENE SUBSTANZEN
C0152426|T019|Q00.1|DMDICD10|CRANIORACHISCHISIS|KRANIORHACHISCHISIS
C0702169|T019|Q00.0|ICD10CM|ANENCEPHALY|ACRANIA
C2879897|T037|T47.92XS|ICD10CM|POISONING BY UNSPECIFIED AGENTS PRIMARILY AFFECTING THE GASTROINTESTINAL SYSTEM, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY UNSP AGENTS AFF THE GI SYS, SELF-HARM, SEQUELA
C2835420|T037|S22.072A|ICD10CM|UNSTABLE BURST FRACTURE OF T9-T10 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSTABLE BURST FRACTURE OF T9-T10 VERTEBRA, INIT FOR CLOS FX
C2835421|T037|S22.072B|ICD10CM|UNSTABLE BURST FRACTURE OF T9-T10 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSTABLE BURST FRACTURE OF T9-T10 VERTEBRA, INIT FOR OPN FX
C2879895|T037|T47.92XA|ICD10CM|POISONING BY UNSPECIFIED AGENTS PRIMARILY AFFECTING THE GASTROINTESTINAL SYSTEM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY UNSP AGENTS AFF THE GI SYS, SELF-HARM, INIT
C0398604|T047|D68.4|ICD10CM|ACQUIRED COAGULATION FACTOR DEFICIENCY|DEFICIENCY OF COAGULATION FACTOR DUE TO LIVER DISEASE
C4237372|T048|F16.959|ICD10CM|HALLUCINOGEN USE, UNSPECIFIED WITH HALLUCINOGEN-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|PHENCYCLIDINE INDUCED PSYCHOTIC DISORDER, WITHOUT USE DISORDER
C2832329|T037|S06.366A|ICD10CM|TRAUMATIC HEMORRHAGE OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|TRAUM HEMOR CEREB, W LOC >24 HR W/O RET CONSC W SURV, INIT
C0042974|T047|D68.0|DMDICD10|VON WILLEBRAND'S DISEASE|WILLEBRAND-JUERGENS-SYNDROM
C0015523|T047|D68.1|DMDICD10|HEREDITARY FACTOR XI DEFICIENCY|HEREDITAERER FAKTOR-XI-MANGEL
C2874715|T048|F16.951|ICD10CM|HALLUCINOGEN USE, UNSPECIFIED WITH HALLUCINOGEN-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|HALLUCINOGEN USE, UNSP W PSYCHOTIC DISORDER W HALLUCINATIONS
C2874714|T048|F16.950|ICD10CM|HALLUCINOGEN USE, UNSPECIFIED WITH HALLUCINOGEN-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|HALLUCINOGEN USE, UNSP W PSYCHOTIC DISORDER W DELUSIONS
C0477316|T047|D68.8|DMDICD10|OTHER SPECIFIED COAGULATION DEFECTS|SONSTIGE NAEHER BEZEICHNETE KOAGULOPATHIEN
C0005779|T047|D68.9|DMDICD10|COAGULATION DEFECT, UNSPECIFIED|KOAGULOPATHIE, NICHT NAEHER BEZEICHNET
C4268399|T047|H40.1114|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, RIGHT EYE, INDETERMINATE STAGE|PRIMARY OPEN-ANGLE GLAUCOMA, RIGHT EYE, INDETERMINATE STAGE
C4268397|T047|H40.1112|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, RIGHT EYE, MODERATE STAGE|PRIMARY OPEN-ANGLE GLAUCOMA, RIGHT EYE, MODERATE STAGE
C4268398|T047|H40.1113|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, RIGHT EYE, SEVERE STAGE|PRIMARY OPEN-ANGLE GLAUCOMA, RIGHT EYE, SEVERE STAGE
C4268395|T047|H40.1110|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, RIGHT EYE, STAGE UNSPECIFIED|PRIMARY OPEN-ANGLE GLAUCOMA, RIGHT EYE, STAGE UNSPECIFIED
C4268396|T047|H40.1111|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, RIGHT EYE, MILD STAGE|PRIMARY OPEN-ANGLE GLAUCOMA, RIGHT EYE, MILD STAGE
C2835327|T037|S22.049B|ICD10CM|UNSPECIFIED FRACTURE OF FOURTH THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF FOURTH THORACIC VERTEBRA, INIT FOR OPN FX
C2835326|T037|S22.049A|ICD10CM|UNSPECIFIED FRACTURE OF FOURTH THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF FOURTH THORACIC VERTEBRA, INIT FOR CLOS FX
C2901416|T046|M84.631A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, RIGHT ULNA, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, RIGHT ULNA, INIT
C2879283|T037|T45.692A|ICD10CM|POISONING BY OTHER FIBRINOLYSIS-AFFECTING DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH FIBRIN-AFFCT DRUGS, SELF-HARM, INIT
C2879285|T037|T45.692S|ICD10CM|POISONING BY OTHER FIBRINOLYSIS-AFFECTING DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH FIBRIN-AFFCT DRUGS, SELF-HARM, SEQUELA
C2896521|T046|M80.029A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, UNSPECIFIED HUMERUS, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, UNSP HUMERUS, INIT
C2833435|T037|S12.390A|ICD10CM|OTHER DISPLACED FRACTURE OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH DISP FX OF FOURTH CERVICAL VERTEBRA, INIT FOR CLOS FX
C2833436|T037|S12.390B|ICD10CM|OTHER DISPLACED FRACTURE OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH DISP FX OF FOURTH CERVICAL VERTEBRA, INIT FOR OPN FX
C4268032|T047|E10.3492|ICD10CM|TYPE 1 DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|TYPE 1 DIAB WITH SEVERE NONP RTNOP WITHOUT MCLR EDEMA, L EYE
C2890304|T037|T83.23XA|ICD10CM|LEAKAGE OF GRAFT OF URINARY ORGAN, INITIAL ENCOUNTER|LEAKAGE OF GRAFT OF URINARY ORGAN, INITIAL ENCOUNTER
C2834066|T037|S14.159S|ICD10CM|OTHER INCOMPLETE LESION AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, SEQUELA|OTH INCMPL LESION AT UNSP LEVEL OF CERV SPINAL CORD, SEQUELA
C2905707|T037|X74.09XA|ICD10CM|INTENTIONAL SELF-HARM BY OTHER GAS, AIR OR SPRING-OPERATED GUN, INITIAL ENCOUNTER|SELF-HARM BY OTH GAS, AIR OR SPRING-OPERATED GUN, INIT
C2858902|T037|S72.464A|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP SUPRCNDL FX W INTRCNDL EXTN LOWER END R FEMUR, INIT
C0349457|T191||ICD10CM|MALIGNANT NEOPLASM OF BODY OF PENIS
C0153599|T191|C60.1|DMDICD10|MALIGNANT NEOPLASM OF GLANS PENIS|BOESARTIGE NEUBILDUNG: GLANS PENIS
C0153598|T191|C60.0|DMDICD10|MALIGNANT NEOPLASM OF PREPUCE|BOESARTIGE NEUBILDUNG: PRAEPUTIUM PENIS
C2834065|T037|S14.159D|ICD10CM|OTHER INCOMPLETE LESION AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|OTH INCMPL LESION AT UNSP LEVEL OF CERV SPINAL CORD, SUBS
C4268809|T046|M84.759A|ICD10CM|COMPLETE OBLIQUE ATYPICAL FEMORAL FRACTURE, UNSPECIFIED LEG, INITIAL ENCOUNTER FOR FRACTURE|COMPLETE OBLIQUE ATYPICAL FEMORAL FRACTURE, UNSP LEG, INIT
C0346225|T191||ICD10CM|MALIGNANT NEOPLASM OF PENIS, UNSPECIFIED
C0349056|T191|C60.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF PENIS|BOESARTIGE NEUBILDUNG: PENIS, MEHRERE TEILBEREICHE UEBERLAPPEND
C2901969|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF LEFT TIBIA
C2901970|T046|M87.063|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED TIBIA|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED TIBIA
C2901968|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF RIGHT TIBIA
C4268118|T047|E11.3593|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|TYPE 2 DIAB WITH PROLIF DIAB RTNOP WITHOUT MACULAR EDEMA, BI
C4268117|T047|E11.3592|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|TYPE 2 DIAB WITH PROLIF DIAB RTNOP WITHOUT MCLR EDEMA, L EYE
C4268116|T047|E11.3591|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|TYPE 2 DIAB WITH PROLIF DIAB RTNOP WITHOUT MCLR EDEMA, R EYE
C2901972|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF LEFT FIBULA
C4509293|T047|L97.305|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED ANKLE WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULCER OF UNSP ANKL WITH MSL INVL W/O EVD OF NECR
C2888680|T047|L97.304|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED ANKLE WITH NECROSIS OF BONE|NON-PRESSURE CHRONIC ULCER OF UNSP ANKLE W NECROSIS OF BONE
C4509294|T047|L97.306|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED ANKLE WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OF UNSP ANKL WITH BONE INVL W/O EVD OF NECR
C2888677|T047|L97.301|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED ANKLE LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHRONIC ULCER OF UNSP ANKLE LIMITED TO BRKDWN SKIN
C4268119|T047|E11.3599|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|TYPE 2 DIAB WITH PROLIF DIAB RTNOP WITHOUT MCLR EDEMA, UNSP
C2888678|T047|L97.302|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED ANKLE WITH FAT LAYER EXPOSED|NON-PRESSURE CHRONIC ULCER OF UNSP ANKLE W FAT LAYER EXPOSED
C2877713|T037|T40.602A|ICD10CM|POISONING BY UNSPECIFIED NARCOTICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY UNSP NARCOTICS, INTENTIONAL SELF-HARM, INIT
C2889345|T047|M05.752|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HIP WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRITIS W RHEU FACTOR OF LEFT HIP W/O ORG/SYS INVOLV
C2889344|T047|M05.751|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT HIP WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRITIS W RHEU FACTOR OF RIGHT HIP W/O ORG/SYS INVOLV
C2896697|T046|M80.829A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, UNSPECIFIED HUMERUS, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, UNSP HUMERUS, INIT
C2832132|T037|S06.319A|ICD10CM|CONTUSION AND LACERATION OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|CONTUS/LAC RIGHT CEREBRUM W LOC OF UNSP DURATION, INIT
C2889346|T047|M05.759|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED HIP WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRITIS W RHEU FACTOR OF UNSP HIP W/O ORG/SYS INVOLV
C2837920|T037|S32.412B|ICD10CM|DISPLACED FRACTURE OF ANTERIOR WALL OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISP FX OF ANTERIOR WALL OF LEFT ACETABULUM, INIT FOR OPN FX
C2900896|T046|M84.422A|ICD10CM|PATHOLOGICAL FRACTURE, LEFT HUMERUS, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, LEFT HUMERUS, INIT FOR FX
C2874582|T048|F14.151|ICD10CM|COCAINE ABUSE WITH COCAINE-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|COCAINE ABUSE W COCAINE-INDUC PSYCHOTIC DISORDER W HALLUCIN
C2874581|T048|F14.150|ICD10CM|COCAINE ABUSE WITH COCAINE-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|COCAINE ABUSE W COCAINE-INDUC PSYCHOTIC DISORDER W DELUSIONS
C0730525|T048||ICD10CM|POST-TRAUMATIC STRESS DISORDER, CHRONIC
C0747767|T048||ICD10CM|POST-TRAUMATIC STRESS DISORDER, ACUTE
C0038436|T048|F43.10|ICD10CM|POST-TRAUMATIC STRESS DISORDER, UNSPECIFIED|POST-TRAUMATIC STRESS DISORDER, UNSPECIFIED
C2882384|T047|I63.419|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF UNSPECIFIED MIDDLE CEREBRAL ARTERY|CEREB INFRC DUE TO EMBOLISM OF UNSP MIDDLE CEREBRAL ARTERY
C2882382|T047|I63.411|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF RIGHT MIDDLE CEREBRAL ARTERY|CEREB INFRC DUE TO EMBOLISM OF RIGHT MIDDLE CEREBRAL ARTERY
C4268485|T047|I63.413|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF BILATERAL MIDDLE CEREBRAL ARTERIES|CEREBRAL INFRC DUE TO EMBOLISM OF BI MIDDLE CEREBRAL ART
C2882383|T047|I63.412|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF LEFT MIDDLE CEREBRAL ARTERY|CEREB INFRC DUE TO EMBOLISM OF LEFT MIDDLE CEREBRAL ARTERY
C2879310|T037|T45.7X2S|ICD10CM|POISONING BY ANTICOAGULANT ANTAGONISTS, VITAMIN K AND OTHER COAGULANTS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY ANTICOAG ANTAG, VIT K AND OTH COAG, SLF-HRM, SQLA
C2857805|T037|S72.326B|ICD10CM|NONDISPLACED TRANSVERSE FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP TRANSVERSE FX SHAFT OF UNSP FEMR, 7THB
C2857806|T037|S72.326C|ICD10CM|NONDISPLACED TRANSVERSE FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP TRANSVERSE FX SHAFT OF UNSP FEMR, 7THC
C2857804|T037|S72.326A|ICD10CM|NONDISPLACED TRANSVERSE FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP TRANSVERSE FRACTURE OF SHAFT OF UNSP FEMUR, INIT
C2874583|T048|F14.159|ICD10CM|COCAINE ABUSE WITH COCAINE-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|COCAINE ABUSE WITH COCAINE-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED
C2858235|T037|S72.391B|ICD10CM|OTHER FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|OTH FX SHAFT OF RIGHT FEMUR, INIT FOR OPN FX TYPE I/2
C2858236|T037|S72.391C|ICD10CM|OTHER FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|OTH FX SHAFT OF RIGHT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2883887|T037|T50.B12A|ICD10CM|POISONING BY SMALLPOX VACCINES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY SMALLPOX VACCINES, INTENTIONAL SELF-HARM, INIT
C2896669|T046|M80.812A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, LEFT SHOULDER, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, L SHOULDER, INIT
C2845970|T191|C79.60|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF UNSPECIFIED OVARY|SECONDARY MALIGNANT NEOPLASM OF UNSPECIFIED OVARY
C1297997|T191|C79.61|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF RIGHT OVARY|SECONDARY MALIGNANT NEOPLASM OF RIGHT OVARY
C1297990|T191|C79.62|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF LEFT OVARY|SECONDARY MALIGNANT NEOPLASM OF LEFT OVARY
C2838607|T037|S34.01XS|ICD10CM|CONCUSSION AND EDEMA OF LUMBAR SPINAL CORD, SEQUELA|CONCUSSION AND EDEMA OF LUMBAR SPINAL CORD, SEQUELA
C2876794|T037|T37.0X2A|ICD10CM|POISONING BY SULFONAMIDES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY SULFONAMIDES, INTENTIONAL SELF-HARM, INIT
C2905666|T037|X71.9XXA|ICD10CM|INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION, UNSPECIFIED, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION, UNSP, INIT
C2838315|T037|S32.482A|ICD10CM|DISPLACED DOME FRACTURE OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED DOME FRACTURE OF LEFT ACETABULUM, INIT FOR CLOS FX
C2838316|T037|S32.482B|ICD10CM|DISPLACED DOME FRACTURE OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISPLACED DOME FRACTURE OF LEFT ACETABULUM, INIT FOR OPN FX
C2838605|T037|S34.01XA|ICD10CM|CONCUSSION AND EDEMA OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|CONCUSSION AND EDEMA OF LUMBAR SPINAL CORD, INIT ENCNTR
C2890686|T037|T84.197A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTERNAL FIXATION DEVICE OF BONE OF LEFT LOWER LEG, INITIAL ENCOUNTER|MECH COMPL OF INT FIX OF BONE OF LEFT LOWER LEG, INIT
C2832694|T037|S06.9X5S|ICD10CM|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, SEQUELA|UNSP INTCRN INJURY W LOC >24 HR W RET CONSC LEV, SEQUELA
C0154754|T047|G60|DMDICD10|HEREDITARY AND IDIOPATHIC NEUROPATHY, UNSPECIFIED|HEREDITAERE UND IDIOPATHISCHE NEUROPATHIE
C2875303|T047|G60.8|ICD10CM|OTHER HEREDITARY AND IDIOPATHIC NEUROPATHIES|RECESSIVELY INHERITED SENSORY NEUROPATHY
C0494493|T047|G60.3|DMDICD10|IDIOPATHIC PROGRESSIVE NEUROPATHY|IDIOPATHISCHE PROGRESSIVE NEUROPATHIE
C0451669|T047|G60.2|DMDICD10|NEUROPATHY IN ASSOCIATION WITH HEREDITARY ATAXIA|NEUROPATHIE IN VERBINDUNG MIT HEREDITAERER ATAXIE
C0282527|T047||ICD10CM|REFSUM'S DISEASE
C2875300|T047|G60.0|ICD10CM|HEREDITARY MOTOR AND SENSORY NEUROPATHY|PERONEAL MUSCULAR ATROPHY (AXONAL TYPE) (HYPERTROPHIC TYPE)
C4270306|T046|T83.491A|ICD10CM|OTHER MECHANICAL COMPLICATION OF IMPLANTED TESTICULAR PROSTHESIS, INITIAL ENCOUNTER|MECH COMPL OF IMPLANTED TESTICULAR PROSTHESIS, INIT
C2712972|T047|K91.850|ICD10CM|POUCHITIS|INFLAMMATION OF INTERNAL ILEOANAL POUCH
C4269410|T037|S02.40ES|ICD10CM|ZYGOMATIC FRACTURE, RIGHT SIDE, SEQUELA|ZYGOMATIC FRACTURE, RIGHT SIDE, SEQUELA
C2833607|T037|S12.631B|ICD10CM|UNSPECIFIED TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP TRAUM NONDISP SPONDYLOLYSIS OF 7TH CERVCAL VERT, 7THB
C2833606|T037|S12.631A|ICD10CM|UNSPECIFIED TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP TRAUM NONDISP SPONDYLOLYSIS OF 7TH CERVCAL VERT, INIT
C2884744|T037|T58.02XS|ICD10CM|TOXIC EFFECT OF CARBON MONOXIDE FROM MOTOR VEHICLE EXHAUST, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFF OF CARB MONX FROM MTR VEH EXHAUST, SLF-HRM, SQLA
C2712860|T046|K91.858|ICD10CM|OTHER COMPLICATIONS OF INTESTINAL POUCH|OTHER COMPLICATIONS OF INTESTINAL POUCH
C2882980|T047|I70.712|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, LEFT LEG|ATHSCL TYPE OF BYPASS OF THE EXTRM W INTRMT CLAUD, LEFT LEG
C2882981|T047|I70.713|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, BILATERAL LEGS|ATHSCL TYPE OF BYPASS OF THE EXTRM W INTRMT CLAUD, BI LEGS
C2874301|T046|E83.30|ICD10CM|DISORDER OF PHOSPHORUS METABOLISM, UNSPECIFIED|DISORDER OF PHOSPHORUS METABOLISM, UNSPECIFIED
C2363067|T047|E83.31|ICD10CM|FAMILIAL HYPOPHOSPHATEMIA|VITAMIN D-RESISTANT OSTEOMALACIA
C2882982|T047|I70.718|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, OTHER EXTREMITY|ATHSCL TYPE OF BYPASS OF THE EXTRM W INTRMT CLAUD, OTH EXTRM
C2882983|T047|I70.719|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, UNSPECIFIED EXTREMITY|ATHSCL TYPE OF BYPASS OF EXTRM W INTRMT CLAUD, UNSP EXTRM
C2856069|T037|S68.626S|ICD10CM|PARTIAL TRAUMATIC TRANSPHALANGEAL AMPUTATION OF RIGHT LITTLE FINGER, SEQUELA|PARTIAL TRAUMATIC TRNSPHAL AMP OF R LITTLE FINGER, SEQUELA
C2888491|T047|L89.504|ICD10CM|PRESSURE ULCER OF UNSPECIFIED ANKLE, STAGE 4|PRESSURE ULCER OF UNSPECIFIED ANKLE, STAGE 4
C2858407|T037|S72.415B|ICD10CM|NONDISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP UNSP CONDYLE FX LOW END L FEMR, 7THB
C2888479|T047|L89.500|ICD10CM|PRESSURE ULCER OF UNSPECIFIED ANKLE, UNSTAGEABLE|PRESSURE ULCER OF UNSPECIFIED ANKLE, UNSTAGEABLE
C2888482|T047|L89.501|ICD10CM|PRESSURE ULCER OF UNSPECIFIED ANKLE, STAGE 1|PRESSURE ULCER OF UNSPECIFIED ANKLE, STAGE 1
C2888485|T047|L89.502|ICD10CM|PRESSURE ULCER OF UNSPECIFIED ANKLE, STAGE 2|PRESSURE ULCER OF UNSPECIFIED ANKLE, STAGE 2
C2888488|T047|L89.503|ICD10CM|PRESSURE ULCER OF UNSPECIFIED ANKLE, STAGE 3|PRESSURE ULCER OF UNSPECIFIED ANKLE, STAGE 3
C2857480|T037|S72.142B|ICD10CM|DISPLACED INTERTROCHANTERIC FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPLACED INTERTROCH FX LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C2857481|T037|S72.142C|ICD10CM|DISPLACED INTERTROCHANTERIC FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPLACED INTERTROCH FX L FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2857479|T037|S72.142A|ICD10CM|DISPLACED INTERTROCHANTERIC FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED INTERTROCHANTERIC FRACTURE OF LEFT FEMUR, INIT
C2888494|T047|L89.509|ICD10CM|PRESSURE ULCER OF UNSPECIFIED ANKLE, UNSPECIFIED STAGE|PRESSURE ULCER OF UNSPECIFIED ANKLE, UNSPECIFIED STAGE
C4270387|T046|T83.718A|ICD10CM|EROSION OF OTHER IMPLANTED MESH TO ORGAN OR TISSUE, INITIAL ENCOUNTER|EROSION OF OTHER IMPLANTED MESH TO ORGAN OR TISSUE, INIT
C2878354|T037|T43.202A|ICD10CM|POISONING BY UNSPECIFIED ANTIDEPRESSANTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY UNSP ANTIDEPRESSANTS, SELF-HARM, INIT
C2853880|T191|C82.99|ICD10CM|FOLLICULAR LYMPHOMA, UNSPECIFIED, EXTRANODAL AND SOLID ORGAN SITES|FOLLICULAR LYMPHOMA, UNSP, EXTRANODAL AND SOLID ORGAN SITES
C2853879|T191|C82.98|ICD10CM|FOLLICULAR LYMPHOMA, UNSPECIFIED, LYMPH NODES OF MULTIPLE SITES|FOLLICULAR LYMPHOMA, UNSP, LYMPH NODES OF MULTIPLE SITES
C2833160|T037|S12.02XB|ICD10CM|UNSTABLE BURST FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSTABLE BURST FX FIRST CERVCAL VERTEBRA, INIT FOR OPN FX
C2833159|T037|S12.02XA|ICD10CM|UNSTABLE BURST FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSTABLE BURST FRACTURE OF FIRST CERVICAL VERTEBRA, INIT
C2853874|T191|C82.93|ICD10CM|FOLLICULAR LYMPHOMA, UNSPECIFIED, INTRA-ABDOMINAL LYMPH NODES|FOLLICULAR LYMPHOMA, UNSP, INTRA-ABDOMINAL LYMPH NODES
C2853873|T191|C82.92|ICD10CM|FOLLICULAR LYMPHOMA, UNSPECIFIED, INTRATHORACIC LYMPH NODES|FOLLICULAR LYMPHOMA, UNSPECIFIED, INTRATHORACIC LYMPH NODES
C2853872|T191|C82.91|ICD10CM|FOLLICULAR LYMPHOMA, UNSPECIFIED, LYMPH NODES OF HEAD, FACE, AND NECK|FOLLICULAR LYMPHOMA, UNSP, NODES OF HEAD, FACE, AND NECK
C2853871|T191|C82.90|ICD10CM|FOLLICULAR LYMPHOMA, UNSPECIFIED, UNSPECIFIED SITE|FOLLICULAR LYMPHOMA, UNSPECIFIED, UNSPECIFIED SITE
C2853878|T191|C82.97|ICD10CM|FOLLICULAR LYMPHOMA, UNSPECIFIED, SPLEEN|FOLLICULAR LYMPHOMA, UNSPECIFIED, SPLEEN
C2853877|T191|C82.96|ICD10CM|FOLLICULAR LYMPHOMA, UNSPECIFIED, INTRAPELVIC LYMPH NODES|FOLLICULAR LYMPHOMA, UNSPECIFIED, INTRAPELVIC LYMPH NODES
C2853876|T191|C82.95|ICD10CM|FOLLICULAR LYMPHOMA, UNSPECIFIED, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|FOLICLAR LYMPHOMA, UNSP, NODES OF ING REGION AND LOWER LIMB
C2853875|T191|C82.94|ICD10CM|FOLLICULAR LYMPHOMA, UNSPECIFIED, LYMPH NODES OF AXILLA AND UPPER LIMB|FOLLICULAR LYMPHOMA, UNSP, NODES OF AXILLA AND UPPER LIMB
C2878072|T037|T42.1X2A|ICD10CM|POISONING BY IMINOSTILBENES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY IMINOSTILBENES, INTENTIONAL SELF-HARM, INIT
C2888844|T047|M00.149|ICD10CM|PNEUMOCOCCAL ARTHRITIS, UNSPECIFIED HAND|PNEUMOCOCCAL ARTHRITIS, UNSPECIFIED HAND
C2854111|T191||ICD10CM|PROLYMPHOCYTIC LEUKEMIA OF T-CELL TYPE, IN RELAPSE
C2869783|T037|S98.111S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT GREAT TOE, SEQUELA|COMPLETE TRAUMATIC AMPUTATION OF RIGHT GREAT TOE, SEQUELA
C2854109|T191|C91.60|ICD10CM|PROLYMPHOCYTIC LEUKEMIA OF T-CELL TYPE NOT HAVING ACHIEVED REMISSION|PROLYMPHOCYTIC LEUKEMIA OF T-CELL TYPE NOT ACHIEVE REMISSION
C2854110|T191||ICD10CM|PROLYMPHOCYTIC LEUKEMIA OF T-CELL TYPE, IN REMISSION
C2888842|T047|M00.141|ICD10CM|PNEUMOCOCCAL ARTHRITIS, RIGHT HAND|PNEUMOCOCCAL ARTHRITIS, RIGHT HAND
C2888843|T047|M00.142|ICD10CM|PNEUMOCOCCAL ARTHRITIS, LEFT HAND|PNEUMOCOCCAL ARTHRITIS, LEFT HAND
C2878074|T037|T42.1X2S|ICD10CM|POISONING BY IMINOSTILBENES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY IMINOSTILBENES, INTENTIONAL SELF-HARM, SEQUELA
C0837750|T047|M08.99|ICD10AM|JUVENILE ARTHRITIS, UNSPECIFIED, MULTIPLE SITES|JUVENILE ARTHRITIS, UNSPECIFIED, SITE UNSPECIFIED
C2889652|T047|M08.98|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, VERTEBRAE|JUVENILE ARTHRITIS, UNSPECIFIED, VERTEBRAE
C2869781|T037|S98.111A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT GREAT TOE, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF RIGHT GREAT TOE, INIT
C2869782|T037|S98.111D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT GREAT TOE, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF RIGHT GREAT TOE, SUBS
C0837750|T047||ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, UNSPECIFIED SITE
C4267892|T047|D89.40|ICD10CM|MAST CELL ACTIVATION, UNSPECIFIED|MAST CELL ACTIVATION DISORDER, UNSPECIFIED
C4267893|T047|D89.41|ICD10CM|MONOCLONAL MAST CELL ACTIVATION SYNDROME|MONOCLONAL MAST CELL ACTIVATION SYNDROME
C4267894|T047|D89.42|ICD10CM|IDIOPATHIC MAST CELL ACTIVATION SYNDROME|IDIOPATHIC MAST CELL ACTIVATION SYNDROME
C4267895|T047|D89.43|ICD10CM|SECONDARY MAST CELL ACTIVATION|SECONDARY MAST CELL ACTIVATION SYNDROME
C3263977|T047|G40.804|ICD10CM|OTHER EPILEPSY, INTRACTABLE, WITHOUT STATUS EPILEPTICUS|OTHER EPILEPSY, INTRACTABLE, WITHOUT STATUS EPILEPTICUS
C3263976|T047|G40.803|ICD10CM|OTHER EPILEPSY, INTRACTABLE, WITH STATUS EPILEPTICUS|OTHER EPILEPSY, INTRACTABLE, WITH STATUS EPILEPTICUS
C4267896|T047|D89.49|ICD10CM|OTHER MAST CELL ACTIVATION DISORDER|OTHER MAST CELL ACTIVATION SYNDROME
C3263973|T047|G40.801|ICD10CM|OTHER EPILEPSY, NOT INTRACTABLE, WITH STATUS EPILEPTICUS|OTHER EPILEPSY WITHOUT INTRACTABILITY WITH STATUS EPILEPTICUS
C2884384|T037|T54.2X2S|ICD10CM|TOXIC EFFECT OF CORROSIVE ACIDS AND ACID-LIKE SUBSTANCES, INTENTIONAL SELF-HARM, SEQUELA|TOX EFF OF CORROSV ACIDS & ACID-LIKE SUBSTNC, SLF-HRM, SQLA
C2901926|T047|M86.652|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, LEFT THIGH|OTHER CHRONIC OSTEOMYELITIS, LEFT THIGH
C2901925|T047|M86.651|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, RIGHT THIGH|OTHER CHRONIC OSTEOMYELITIS, RIGHT THIGH
C2901927|T047|M86.65|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, UNSPECIFIED THIGH|OTHER CHRONIC OSTEOMYELITIS, THIGH
C2884382|T037|T54.2X2A|ICD10CM|TOXIC EFFECT OF CORROSIVE ACIDS AND ACID-LIKE SUBSTANCES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOX EFF OF CORROSV ACIDS & ACID-LIKE SUBSTNC, SLF-HRM, INIT
C2887933|T047|K72.01|ICD10CM|ACUTE AND SUBACUTE HEPATIC FAILURE WITH COMA|ACUTE AND SUBACUTE HEPATIC FAILURE WITH COMA
C1406683|T047||ICD10CM|POSTSURGICAL MALABSORPTION, NOT ELSEWHERE CLASSIFIED
C2842097|T191|C50.229|ICD10CM|MALIGNANT NEOPLASM OF UPPER-INNER QUADRANT OF UNSPECIFIED MALE BREAST|MALIG NEOPLASM OF UPPER-INNER QUADRANT OF UNSP MALE BREAST
C2842096|T191|C50.222|ICD10CM|MALIGNANT NEOPLASM OF UPPER-INNER QUADRANT OF LEFT MALE BREAST|MALIG NEOPLASM OF UPPER-INNER QUADRANT OF LEFT MALE BREAST
C2842095|T191|C50.221|ICD10CM|MALIGNANT NEOPLASM OF UPPER-INNER QUADRANT OF RIGHT MALE BREAST|MALIG NEOPLASM OF UPPER-INNER QUADRANT OF RIGHT MALE BREAST
C2874023|T047|E10.21|ICD10CM|TYPE 1 DIABETES MELLITUS WITH DIABETIC NEPHROPATHY|TYPE 1 DIABETES MELLITUS WITH INTRACAPILLARY GLOMERULONEPHROSIS
C0432429|T047|Q92.1|DMDICD10|WHOLE CHROMOSOME TRISOMY, MOSAICISM (MITOTIC NONDISJUNCTION)|VOLLSTAENDIGE TRISOMIE, MOSAIK (MITOTISCHE NON-DISJUNCTION)
C2910358|T019|Q92.2|ICD10CM|PARTIAL TRISOMY|WHOLE ARM OR MORE DUPLICATED
C2874025|T047|E10.22|ICD10CM|TYPE 1 DIABETES MELLITUS WITH DIABETIC CHRONIC KIDNEY DISEASE|TYPE 1 DIABETES MELLITUS W DIABETIC CHRONIC KIDNEY DISEASE
C2910359|T047|Q92.5|ICD10CM|DUPLICATIONS WITH OTHER COMPLEX REARRANGEMENTS|PARTIAL TRISOMY DUE TO UNBALANCED TRANSLOCATIONS
C0432435|T049|Q92.7|DMDICD10|TRIPLOIDY AND POLYPLOIDY|TRIPLOIDIE UND POLYPLOIDIE
C2874027|T047|E10.29|ICD10CM|TYPE 1 DIABETES MELLITUS WITH OTHER DIABETIC KIDNEY COMPLICATION|TYPE 1 DIABETES MELLITUS W OTH DIABETIC KIDNEY COMPLICATION
C0495649|T047|Q92.9|DMDICD10|TRISOMY AND PARTIAL TRISOMY OF AUTOSOMES, UNSPECIFIED|TRISOMIE UND PARTIELLE TRISOMIE DER AUTOSOMEN, NICHT NAEHER BEZEICHNET
C2832477|T037|S06.5X2A|ICD10CM|TRAUMATIC SUBDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|TRAUM SUBDR HEM W LOSS OF CONSCIOUSNESS OF 31-59 MIN, INIT
C2832479|T037|S06.5X2S|ICD10CM|TRAUMATIC SUBDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|TRAUM SUBDR HEM W LOC OF 31-59 MIN, SEQUELA
C2889244|T047|M05.439|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSP WRIST
C4268007|T047|E09.37X1|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, RIGHT EYE|DRUG/CHEM DIAB W DIAB MCLR EDMA, RESOLVED FOL TRTMT, R EYE
C4268009|T047|E09.37X3|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, BILATERAL|DRUG/CHEM DIAB WITH DIAB MCLR EDEMA, RESOLVED FOL TRTMT, BI
C4268008|T047|E09.37X2|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, LEFT EYE|DRUG/CHEM DIAB W DIAB MCLR EDMA, RESOLVED FOL TRTMT, L EYE
C2889243|T047|M05.432|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT WRIST|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889242|T047|M05.431|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT WRIST|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT WRIST
C4268010|T047|E09.37X9|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, UNSPECIFIED EYE|DRUG/CHEM DIAB WITH DIAB MCLR EDMA, RESOLVED FOL TRTMT, UNSP
C2874277|T047|E76.210|ICD10CM|MORQUIO A MUCOPOLYSACCHARIDOSES|MORQUIO A MUCOPOLYSACCHARIDOSES
C0349074|T046|I23.4|DMDICD10|RUPTURE OF CHORDAE TENDINEAE AS CURRENT COMPLICATION FOLLOWING ACUTE MYOCARDIAL INFARCTION|RUPTUR DER CHORDAE TENDINEAE ALS AKUTE KOMPLIKATION NACH AKUTEM MYOKARDINFARKT
C3665604|T047|I23.5|DMDICD10|RUPTURE OF PAPILLARY MUSCLE AS CURRENT COMPLICATION FOLLOWING ACUTE MYOCARDIAL INFARCTION|PAPILLARMUSKELRUPTUR ALS AKUTE KOMPLIKATION NACH AKUTEM MYOKARDINFARKT
C2878328|T037|T43.1X2A|ICD10CM|POISONING BY MONOAMINE-OXIDASE-INHIBITOR ANTIDEPRESSANTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY MAO INHIB ANTIDEPRESSANTS, SELF-HARM, INIT
C2901408|T046|M84.629A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, UNSPECIFIED HUMERUS, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, UNSP HUMERUS, INIT
C0348876|T047|I23.6|DMDICD10|THROMBOSIS OF ATRIUM, AURICULAR APPENDAGE, AND VENTRICLE AS CURRENT COMPLICATIONS FOLLOWING ACUTE MYOCARDIAL INFARCTION|THROMBOSE DES VORHOFES, DES HERZOHRES ODER DER KAMMER ALS AKUTE KOMPLIKATION NACH AKUTEM MYOKARDINFARKT
C2835754|T037|S24.0XXS|ICD10CM|CONCUSSION AND EDEMA OF THORACIC SPINAL CORD, SEQUELA|CONCUSSION AND EDEMA OF THORACIC SPINAL CORD, SEQUELA
C2879207|T037|T45.602S|ICD10CM|POISONING BY UNSPECIFIED FIBRINOLYSIS-AFFECTING DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY UNSP FIBRIN-AFFCT DRUGS, SELF-HARM, SEQUELA
C0494662|T047|J61|DMDICD10|PNEUMOCONIOSIS DUE TO ASBESTOS AND OTHER MINERAL FIBERS|PNEUMOKONIOSE DURCH ASBEST UND SONSTIGE ANORGANISCHE FASERN
C0003165|T047|J60|DMDICD10|COALWORKER'S PNEUMOCONIOSIS|KOHLENBERGARBEITER-PNEUMOKONIOSE
C2887470|T047|J65|ICD10CM|PNEUMOCONIOSIS ASSOCIATED WITH TUBERCULOSIS|ANY CONDITION IN J60-J64 WITH TUBERCULOSIS, ANY TYPE IN A15
C0032273|T047|J64|DMDICD10|UNSPECIFIED PNEUMOCONIOSIS|NICHT NAEHER BEZEICHNETE PNEUMOKONIOSE
C2835752|T037|S24.0XXA|ICD10CM|CONCUSSION AND EDEMA OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|CONCUSSION AND EDEMA OF THORACIC SPINAL CORD, INIT ENCNTR
C2901474|T046|M84.650A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, PELVIS, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, PELVIS, INIT FOR FX
C2835753|T037|S24.0XXD|ICD10CM|CONCUSSION AND EDEMA OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|CONCUSSION AND EDEMA OF THORACIC SPINAL CORD, SUBS ENCNTR
C2879205|T037|T45.602A|ICD10CM|POISONING BY UNSPECIFIED FIBRINOLYSIS-AFFECTING DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY UNSP FIBRIN-AFFCT DRUGS, SELF-HARM, INIT
C4270299|T046|T83.421A|ICD10CM|DISPLACEMENT OF IMPLANTED TESTICULAR PROSTHESIS, INITIAL ENCOUNTER|DISPLACEMENT OF IMPLANTED TESTICULAR PROSTHESIS, INIT
C2858509|T037|S72.425B|ICD10CM|NONDISPLACED FRACTURE OF LATERAL CONDYLE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF LATERAL CONDYLE OF L FEMR, 7THB
C2858510|T037|S72.425C|ICD10CM|NONDISPLACED FRACTURE OF LATERAL CONDYLE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF LATERAL CONDYLE OF L FEMR, 7THC
C2858508|T037|S72.425A|ICD10CM|NONDISPLACED FRACTURE OF LATERAL CONDYLE OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF LATERAL CONDYLE OF LEFT FEMUR, INIT
C2832429|T037|S06.4X0A|ICD10CM|EPIDURAL HEMORRHAGE WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|EPIDURAL HEMORRHAGE W/O LOSS OF CONSCIOUSNESS, INIT ENCNTR
C2830423|T033|R40.2340|ICD10CM|COMA SCALE, BEST MOTOR RESPONSE, FLEXION WITHDRAWAL, UNSPECIFIED TIME|COMA SCALE, BEST MOTOR, FLEXION WITHDRAWAL, UNSP TIME
C2830424|T033|R40.2341|ICD10CM|COMA SCALE, BEST MOTOR RESPONSE, FLEXION WITHDRAWAL, IN THE FIELD [EMT OR AMBULANCE]|COMA SCALE, BEST MOTOR, FLEXION WITHDRAWAL, IN THE FIELD
C2830425|T033|R40.2342|ICD10CM|COMA SCALE, BEST MOTOR RESPONSE, FLEXION WITHDRAWAL, AT ARRIVAL TO EMERGENCY DEPARTMENT|COMA SCALE, BEST MOTOR RESPONSE, FLEXION WITHDRAWAL, EMR
C2830426|T033|R40.2343|ICD10CM|COMA SCALE, BEST MOTOR RESPONSE, FLEXION WITHDRAWAL, AT HOSPITAL ADMISSION|COMA SCALE, BEST MOTOR RESPONSE, FLEXION WITHDRAWAL, ADMIT
C2830427|T033|R40.2344|ICD10CM|COMA SCALE, BEST MOTOR RESPONSE, FLEXION WITHDRAWAL, 24 HOURS OR MORE AFTER HOSPITAL ADMISSION|COMA SCALE, BEST MOTOR RESPONSE, FLEXION WITHDRAWAL, 24+HRS
C2832439|T037|S06.4X2S|ICD10CM|EPIDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|EPIDURAL HEMORRHAGE W LOC OF 31-59 MIN, SEQUELA
C2832437|T037|S06.4X2A|ICD10CM|EPIDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|EPIDURAL HEMORRHAGE W LOC OF 31-59 MIN, INIT
C2855889|T037|S68.116S|ICD10CM|COMPLETE TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF RIGHT LITTLE FINGER, SEQUELA|COMPLETE TRAUMATIC MCP AMP OF R LITTLE FINGER, SEQUELA
C2878281|T037|T43.012S|ICD10CM|POISONING BY TRICYCLIC ANTIDEPRESSANTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY TRICYCLIC ANTIDEPRESSANTS, SELF-HARM, SEQUELA
C0343491|T047|A39.84|ICD10CM|POSTMENINGOCOCCAL ARTHRITIS|POSTMENINGOCOCCAL ARTHRITIS
C2878279|T037|T43.012A|ICD10CM|POISONING BY TRICYCLIC ANTIDEPRESSANTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY TRICYCLIC ANTIDEPRESSANTS, SELF-HARM, INIT
C2856501|T037|S72.002C|ICD10CM|FRACTURE OF UNSPECIFIED PART OF NECK OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|FX UNSP PART OF NECK OF L FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C1457881|T047|A39.83|ICD10CM|MENINGOCOCCAL ARTHRITIS|MENINGOCOCCAL ARTHRITIS
C2902036|T046|M87.219|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED SHOULDER|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED SHOULDER
C2891331|T046||ICD10CM|INFECTION OF AMPUTATION STUMP, LEFT UPPER EXTREMITY
C2856500|T037|S72.002B|ICD10CM|FRACTURE OF UNSPECIFIED PART OF NECK OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|FX UNSP PART OF NECK OF LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C2902034|T046|M87.211|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, RIGHT SHOULDER|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, RIGHT SHOULDER
C2884464|T037|T56.0X2A|ICD10CM|TOXIC EFFECT OF LEAD AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF LEAD AND ITS COMPOUNDS, SELF-HARM, INIT
C2902035|T046|M87.212|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, LEFT SHOULDER|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, LEFT SHOULDER
C2882075|T047|I11.9|ICD10CM|HYPERTENSIVE HEART DISEASE WITHOUT HEART FAILURE|HYPERTENSIVE HEART DISEASE WITHOUT HEART FAILURE
C2889435|T047|M06.271|ICD10CM|RHEUMATOID BURSITIS, RIGHT ANKLE AND FOOT|RHEUMATOID BURSITIS, RIGHT ANKLE AND FOOT
C2889436|T047|M06.272|ICD10CM|RHEUMATOID BURSITIS, LEFT ANKLE AND FOOT|RHEUMATOID BURSITIS, LEFT ANKLE AND FOOT
C1400066|T047|I11.0|ICD10CM|HYPERTENSIVE HEART DISEASE WITH HEART FAILURE|HYPERTENSIVE HEART DISEASE WITH HEART FAILURE
C4269420|T037|S02.600B|ICD10CM|FRACTURE OF UNSPECIFIED PART OF BODY OF MANDIBLE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FX UNSP PART OF BODY OF MANDIBLE, UNSPECIFIED SIDE, 7THB
C2884466|T037|T56.0X2S|ICD10CM|TOXIC EFFECT OF LEAD AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF LEAD AND ITS COMPOUNDS, SELF-HARM, SEQUELA
C2889437|T047|M06.279|ICD10CM|RHEUMATOID BURSITIS, UNSPECIFIED ANKLE AND FOOT|RHEUMATOID BURSITIS, UNSPECIFIED ANKLE AND FOOT
C2891332|T046||ICD10CM|INFECTION OF AMPUTATION STUMP, RIGHT LOWER EXTREMITY
C2888031|T046|K94.30|ICD10CM|ESOPHAGOSTOMY COMPLICATIONS, UNSPECIFIED|ESOPHAGOSTOMY COMPLICATIONS, UNSPECIFIED
C2888032|T046|K94.31|ICD10CM|ESOPHAGOSTOMY HEMORRHAGE|ESOPHAGOSTOMY HEMORRHAGE
C1456233|T046|K94.32|ICD10CM|ESOPHAGOSTOMY INFECTION|ESOPHAGOSTOMY INFECTION
C1456235|T046|K94.33|ICD10CM|ESOPHAGOSTOMY MALFUNCTION|ESOPHAGOSTOMY MALFUNCTION
C2888033|T047|K94.39|ICD10CM|OTHER COMPLICATIONS OF ESOPHAGOSTOMY|OTHER COMPLICATIONS OF ESOPHAGOSTOMY
C2879442|T037|T46.2X2S|ICD10CM|POISONING BY OTHER ANTIDYSRHYTHMIC DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH ANTIDYSRHYTHMIC DRUGS, SELF-HARM, SEQUELA
C2880106|T047|A06.5|ICD10CM|AMEBIC LUNG ABSCESS|AMEBIC ABSCESS OF LUNG (AND LIVER)
C2837839|T037|S32.313A|ICD10CM|DISPLACED AVULSION FRACTURE OF UNSPECIFIED ILIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED AVULSION FRACTURE OF UNSP ILIUM, INIT FOR CLOS FX
C2889442|T046|M06.319|ICD10CM|RHEUMATOID NODULE, UNSPECIFIED SHOULDER|RHEUMATOID NODULE, UNSPECIFIED SHOULDER
C2889441|T046|M06.312|ICD10CM|RHEUMATOID NODULE, LEFT SHOULDER|RHEUMATOID NODULE, LEFT SHOULDER
C2889440|T046|M06.311|ICD10CM|RHEUMATOID NODULE, RIGHT SHOULDER|RHEUMATOID NODULE, RIGHT SHOULDER
C2891330|T046||ICD10CM|INFECTION OF AMPUTATION STUMP, RIGHT UPPER EXTREMITY
C0153405|T191|C14.0|DMDICD10|MALIGNANT NEOPLASM OF PHARYNX, UNSPECIFIED|BOESARTIGE NEUBILDUNG: PHARYNX, NICHT NAEHER BEZEICHNET
C2885239|T037|T62.1X2S|ICD10CM|TOXIC EFFECT OF INGESTED BERRIES, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF INGESTED BERRIES, SELF-HARM, SEQUELA
C0153516|T191|C41.4|DMDICD10|MALIGNANT NEOPLASM OF PELVIC BONES, SACRUM AND COCCYX|BOESARTIGE NEUBILDUNG DES KNOCHENS UND DES GELENKKNORPELS: BECKENKNOCHEN
C0346667|T191|C41.2|DMDICD10|MALIGNANT NEOPLASM OF VERTEBRAL COLUMN|BOESARTIGE NEUBILDUNG DES KNOCHENS UND DES GELENKKNORPELS: WIRBELSAEULE
C0153513|T191|C41.3|DMDICD10|MALIGNANT NEOPLASM OF RIBS, STERNUM AND CLAVICLE|BOESARTIGE NEUBILDUNG DES KNOCHENS UND DES GELENKKNORPELS: RIPPEN, STERNUM UND KLAVIKULA
C0346665|T191|C41.0|ICD10CM|MALIGNANT NEOPLASM OF BONES OF SKULL AND FACE|MALIGNANT NEOPLASM OF MAXILLA (SUPERIOR)
C0153511|T191|C41.1|DMDICD10|MALIGNANT NEOPLASM OF MANDIBLE|BOESARTIGE NEUBILDUNG DES KNOCHENS UND DES GELENKKNORPELS: UNTERKIEFERKNOCHEN
C2837931|T191|C14.8|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF LIP, ORAL CAVITY AND PHARYNX|PRIMARY MALIGNANT NEOPLASM OF TWO OR MORE CONTIGUOUS SITES OF LIP, ORAL CAVITY AND PHARYNX
C2896492|T046|M80.012A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, LEFT SHOULDER, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, L SHOULDER, INIT
C0153509|T191|C41.9|DMDICD10|MALIGNANT NEOPLASM OF BONE AND ARTICULAR CARTILAGE, UNSPECIFIED|BOESARTIGE NEUBILDUNG: KNOCHEN UND GELENKKNORPEL, NICHT NAEHER BEZEICHNET
C2888645|T047|L97.111|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT THIGH LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHRONIC ULCER OF RIGHT THIGH LIMITED TO BRKDWN SKIN
C2888646|T047|L97.112|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT THIGH WITH FAT LAYER EXPOSED|NON-PRS CHRONIC ULCER OF RIGHT THIGH W FAT LAYER EXPOSED
C2888647|T047|L97.113|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT THIGH WITH NECROSIS OF MUSCLE|NON-PRS CHRONIC ULCER OF RIGHT THIGH W NECROSIS OF MUSCLE
C2888648|T047|L97.114|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT THIGH WITH NECROSIS OF BONE|NON-PRESSURE CHRONIC ULCER OF RIGHT THIGH W NECROSIS OF BONE
C4509278|T047|L97.115|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT THIGH WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULCER OF R THIGH WITH MSL INVL W/O EVD OF NECR
C4509279|T047|L97.116|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT THIGH WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULCER OF R THIGH WITH BONE INVL W/O EVD OF NECR
C2835811|T037|S24.134S|ICD10CM|ANTERIOR CORD SYNDROME AT T11-T12 LEVEL OF THORACIC SPINAL CORD, SEQUELA|ANTERIOR CORD SYNDROME AT T11-T12, SEQUELA
C4509280|T047|L97.118|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT THIGH WITH OTHER SPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF RIGHT THIGH WITH OTH SEVERITY
C2888649|T047|L97.119|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT THIGH WITH UNSPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF RIGHT THIGH WITH UNSP SEVERITY
C2861668|T191|D03.20|ICD10CM|MELANOMA IN SITU OF UNSPECIFIED EAR AND EXTERNAL AURICULAR CANAL|MELANOMA IN SITU OF UNSP EAR AND EXTERNAL AURICULAR CANAL
C2837956|T191|C34.32|ICD10CM|MALIGNANT NEOPLASM OF LOWER LOBE, LEFT BRONCHUS OR LUNG|MALIGNANT NEOPLASM OF LOWER LOBE, LEFT BRONCHUS OR LUNG
C2861670|T191|D03.22|ICD10CM|MELANOMA IN SITU OF LEFT EAR AND EXTERNAL AURICULAR CANAL|MELANOMA IN SITU OF LEFT EAR AND EXTERNAL AURICULAR CANAL
C2845902|T191|C69.10|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED CORNEA|MALIGNANT NEOPLASM OF UNSPECIFIED CORNEA
C2885253|T037|T62.2X2A|ICD10CM|TOXIC EFFECT OF OTHER INGESTED (PARTS OF) PLANT(S), INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF INGESTED (PARTS OF) PLANT(S), SLF-HRM, INIT
C2837955|T191|C34.31|ICD10CM|MALIGNANT NEOPLASM OF LOWER LOBE, RIGHT BRONCHUS OR LUNG|MALIGNANT NEOPLASM OF LOWER LOBE, RIGHT BRONCHUS OR LUNG
C2902914|T047|N06.8|ICD10CM|ISOLATED PROTEINURIA WITH OTHER MORPHOLOGIC LESION|ISOLATED PROTEINURIA WITH OTHER MORPHOLOGIC LESION
C2902915|T047|N06.9|ICD10CM|ISOLATED PROTEINURIA WITH UNSPECIFIED MORPHOLOGIC LESION|ISOLATED PROTEINURIA WITH UNSPECIFIED MORPHOLOGIC LESION
C0495040|T047|N06.4|DMDICD10|ISOLATED PROTEINURIA WITH DIFFUSE ENDOCAPILLARY PROLIFERATIVE GLOMERULONEPHRITIS|ISOLIERTE PROTEINURIE MIT ANGABE MORPHOLOGISCHER VERAENDERUNGEN: DIFFUSE ENDOKAPILLAER-PROLIFERATIVE GLOMERULONEPHRITIS
C2902910|T033|N06.5|ICD10CM|ISOLATED PROTEINURIA WITH DIFFUSE MESANGIOCAPILLARY GLOMERULONEPHRITIS|ISOLATED PROTEINURIA WITH MEMBRANOPROLIFERATIVE GLOMERULONEPHRITIS, TYPES 1 AND 3, OR NOS
C2902911|T033|N06.6|ICD10CM|ISOLATED PROTEINURIA WITH DENSE DEPOSIT DISEASE|ISOLATED PROTEINURIA WITH MEMBRANOPROLIFERATIVE GLOMERULONEPHRITIS, TYPE 2
C2902912|T033|N06.7|ICD10CM|ISOLATED PROTEINURIA WITH DIFFUSE CRESCENTIC GLOMERULONEPHRITIS|ISOLATED PROTEINURIA WITH EXTRACAPILLARY GLOMERULONEPHRITIS
C2902906|T033|N06.0|ICD10CM|ISOLATED PROTEINURIA WITH MINOR GLOMERULAR ABNORMALITY|ISOLATED PROTEINURIA WITH MINIMAL CHANGE LESION
C2902909|T033|N06.1|ICD10CM|ISOLATED PROTEINURIA WITH FOCAL AND SEGMENTAL GLOMERULAR LESIONS|ISOLATED PROTEINURIA WITH FOCAL GLOMERULONEPHRITIS
C0495038|T047|N06.2|DMDICD10|ISOLATED PROTEINURIA WITH DIFFUSE MEMBRANOUS GLOMERULONEPHRITIS|ISOLIERTE PROTEINURIE MIT ANGABE MORPHOLOGISCHER VERAENDERUNGEN: DIFFUSE MEMBRANOESE GLOMERULONEPHRITIS
C0495039|T047|N06.3|DMDICD10|ISOLATED PROTEINURIA WITH DIFFUSE MESANGIAL PROLIFERATIVE GLOMERULONEPHRITIS|ISOLIERTE PROTEINURIE MIT ANGABE MORPHOLOGISCHER VERAENDERUNGEN: DIFFUSE MESANGIOPROLIFERATIVE GLOMERULONEPHRITIS
C0342844|T047|E77|DMDICD10|DISORDER OF GLYCOPROTEIN METABOLISM, UNSPECIFIED|STOERUNGEN DES GLYKOPROTEINSTOFFWECHSELS
C0348493|T047|E77.8|DMDICD10|OTHER DISORDERS OF GLYCOPROTEIN METABOLISM|SONSTIGE STOERUNGEN DES GLYKOPROTEINSTOFFWECHSELS
C2838393|T037|S32.519A|ICD10CM|FRACTURE OF SUPERIOR RIM OF UNSPECIFIED PUBIS, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF SUPERIOR RIM OF UNSP PUBIS, INIT FOR CLOS FX
C1257960|T047|E77.1|ICD10CM|DEFECTS IN GLYCOPROTEIN DEGRADATION|MANNOSIDOSIS
C2874286|T047|E77.0|ICD10CM|DEFECTS IN POST-TRANSLATIONAL MODIFICATION OF LYSOSOMAL ENZYMES|MUCOLIPIDOSIS III [PSEUDO-HURLER POLYDYSTROPHY]
C2891333|T046||ICD10CM|INFECTION OF AMPUTATION STUMP, LEFT LOWER EXTREMITY
C2877946|T037|T41.292A|ICD10CM|POISONING BY OTHER GENERAL ANESTHETICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH GENERAL ANESTHETICS, SELF-HARM, INIT
C4267874|T191|C81.76|ICD10CM|OTHER HODGKIN LYMPHOMA, INTRAPELVIC LYMPH NODES|OTHER HODGKIN LYMPHOMA, INTRAPELVIC LYMPH NODES
C4267875|T191|C81.77|ICD10CM|OTHER HODGKIN LYMPHOMA, SPLEEN|OTHER HODGKIN LYMPHOMA, SPLEEN
C4267872|T191|C81.74|ICD10CM|OTHER HODGKIN LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB|OTHER HODGKIN LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB
C4267873|T191|C81.75|ICD10CM|OTHER HODGKIN LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|OTHER HODGKIN LYMPHOMA, NODES OF ING REGION AND LOWER LIMB
C4267870|T191|C81.72|ICD10CM|OTHER HODGKIN LYMPHOMA, INTRATHORACIC LYMPH NODES|OTHER HODGKIN LYMPHOMA, INTRATHORACIC LYMPH NODES
C4267871|T191|C81.73|ICD10CM|OTHER HODGKIN LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES|OTHER HODGKIN LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES
C4267868|T191|C81.70|ICD10CM|OTHER HODGKIN LYMPHOMA, UNSPECIFIED SITE|OTHER HODGKIN LYMPHOMA, UNSPECIFIED SITE
C4267869|T191|C81.71|ICD10CM|OTHER HODGKIN LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK|OTHER HODGKIN LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK
C4267876|T191|C81.78|ICD10CM|OTHER HODGKIN LYMPHOMA, LYMPH NODES OF MULTIPLE SITES|OTHER HODGKIN LYMPHOMA, LYMPH NODES OF MULTIPLE SITES
C4267877|T191|C81.79|ICD10CM|OTHER HODGKIN LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES|OTHER HODGKIN LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES
C0343539|T047|A81.8|ICD10CM|OTHER ATYPICAL VIRUS INFECTIONS OF CENTRAL NERVOUS SYSTEM|OTHER ATYPICAL VIRUS INFECTIONS OF CENTRAL NERVOUS SYSTEM
C0022802|T047|A81.81|ICD10CM|KURU|KURU
C0206042|T047|A81.83|ICD10CM|FATAL FAMILIAL INSOMNIA|FFI
C0017495|T047|A81.82|ICD10CM|GERSTMANN-STRAUSSLER-SCHEINKER SYNDROME|GSS SYNDROME
C2889015|T046|M02.169|ICD10CM|POSTDYSENTERIC ARTHROPATHY, UNSPECIFIED KNEE|POSTDYSENTERIC ARTHROPATHY, UNSPECIFIED KNEE
C2832370|T037|S06.376A|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF CEREBELLUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|CONTUS/LAC/HEM CRBLM W LOC >24 HR W/O RET CONSC W SURV, INIT
C2886176|T037|T65.832A|ICD10CM|TOXIC EFFECT OF FIBERGLASS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF FIBERGLASS, INTENTIONAL SELF-HARM, INIT
C2889013|T047|M02.161|ICD10CM|POSTDYSENTERIC ARTHROPATHY, RIGHT KNEE|POSTDYSENTERIC ARTHROPATHY, RIGHT KNEE
C2889014|T047|M02.162|ICD10CM|POSTDYSENTERIC ARTHROPATHY, LEFT KNEE|POSTDYSENTERIC ARTHROPATHY, LEFT KNEE
C2889396|T047|M06.03|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, UNSPECIFIED WRIST|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, WRIST
C0840029|T046|M87.29|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, MULTIPLE SITES|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, MULTIPLE SITES
C2901162|T046|M84.521A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, RIGHT HUMERUS, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, R HUMERUS, INIT
C2901335|T046|M84.574A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, RIGHT FOOT, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, RIGHT FOOT, INIT
C2901184|T046|M84.531A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, RIGHT ULNA, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, RIGHT ULNA, INIT
C2886178|T037|T65.832S|ICD10CM|TOXIC EFFECT OF FIBERGLASS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF FIBERGLASS, INTENTIONAL SELF-HARM, SEQUELA
C2887193|T047|I83.024|ICD10CM|VARICOSE VEINS OF LEFT LOWER EXTREMITY WITH ULCER OF HEEL AND MIDFOOT|VARICOSE VEINS OF L LOW EXTREM W ULCER OF HEEL AND MIDFOOT
C2874472|T048||ICD10CM|CANNABIS ABUSE WITH INTOXICATION, UNCOMPLICATED
C2874473|T048|F12.121|ICD10CM|CANNABIS ABUSE WITH INTOXICATION DELIRIUM|CANNABIS ABUSE WITH INTOXICATION DELIRIUM
C2874474|T048|F12.122|ICD10CM|CANNABIS ABUSE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE|CANNABIS ABUSE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE
C4268225|T048|F13.24|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED MOOD DISORDER|SEDATIVE, HYPNOTIC, OR ANXIOLYTIC USE DISORDER, SEVERE, WITH SEDATIVE, HYPNOTIC, OR ANXIOLYTIC-INDUCED DEPRESSIVE DISORDER
C4268227|T048|F13.27|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED PERSISTING DEMENTIA|SEDATIVE, HYPNOTIC, OR ANXIOLYTIC USE DISORDER, SEVERE, WITH SEDATIVE, HYPNOTIC, OR ANXIOLYTIC-INDUCED MAJOR NEUROCOGNITIVE DISORDER
C2874543|T048|F13.26|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED PERSISTING AMNESTIC DISORDER|SEDATV/HYP/ANXIOLYTC DEPEND W PERSISTING AMNESTIC DISORDER
C2874549|T048|F13.29|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH UNSPECIFIED SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED DISORDER|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE W UNSP DISORDER
C2874475|T048|F12.129|ICD10CM|CANNABIS ABUSE WITH INTOXICATION, UNSPECIFIED|CANNABIS ABUSE WITH INTOXICATION, UNSPECIFIED
C2873870|T047|E05.21|ICD10CM|THYROTOXICOSIS WITH TOXIC MULTINODULAR GOITER WITH THYROTOXIC CRISIS OR STORM|THYROTXCOSIS W TOXIC MULTINODULAR GOITER W THYROTOXIC CRISIS
C2873869|T047|E05.20|ICD10CM|THYROTOXICOSIS WITH TOXIC MULTINODULAR GOITER WITHOUT THYROTOXIC CRISIS OR STORM|THYROTXCOSIS W TOXIC MULTINOD GOITER W/O THYROTOXIC CRISIS
C4269312|T037|S02.11ES|ICD10CM|TYPE III OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, SEQUELA|TYPE III OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, SEQUELA
C2905769|T037|X79.XXXA|ICD10CM|INTENTIONAL SELF-HARM BY BLUNT OBJECT, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY BLUNT OBJECT, INITIAL ENCOUNTER
C4269308|T037|S02.11EB|ICD10CM|TYPE III OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE III OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, 7THB
C4269307|T037|S02.11EA|ICD10CM|TYPE III OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE III OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, INIT
C2905770|T037|X79.XXXD|ICD10CM|INTENTIONAL SELF-HARM BY BLUNT OBJECT, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY BLUNT OBJECT, SUBSEQUENT ENCOUNTER
C2833450|T037|S12.400A|ICD10CM|UNSPECIFIED DISPLACED FRACTURE OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP DISP FX OF FIFTH CERVICAL VERTEBRA, INIT FOR CLOS FX
C2833451|T037|S12.400B|ICD10CM|UNSPECIFIED DISPLACED FRACTURE OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP DISP FX OF FIFTH CERVICAL VERTEBRA, INIT FOR OPN FX
C3263939|T191|C93.Z0|ICD10CM|OTHER MONOCYTIC LEUKEMIA, NOT HAVING ACHIEVED REMISSION|OTHER MONOCYTIC LEUKEMIA, NOT HAVING ACHIEVED REMISSION
C0153905|T191|C93.Z1|ICD10CM|OTHER MONOCYTIC LEUKEMIA, IN REMISSION|OTHER MONOCYTIC LEUKEMIA, IN REMISSION
C2349293|T191|C93.Z2|ICD10CM|OTHER MONOCYTIC LEUKEMIA, IN RELAPSE|OTHER MONOCYTIC LEUKEMIA, IN RELAPSE
C2901899|T047|M86.539|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED RADIUS AND ULNA|OTH CHRONIC HEMATOGENOUS OSTEOMYELITIS, UNSP RADIUS AND ULNA
C2901898|T047|M86.532|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, LEFT RADIUS AND ULNA|OTH CHRONIC HEMATOGENOUS OSTEOMYELITIS, LEFT RADIUS AND ULNA
C2901897|T047|M86.531|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, RIGHT RADIUS AND ULNA|OTH CHRONIC HEMATOGENOUS OSTEOMYELIT, RIGHT RADIUS AND ULNA
C2857445|T037|S72.136A|ICD10CM|NONDISPLACED APOPHYSEAL FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED APOPHYSEAL FRACTURE OF UNSP FEMUR, INIT
C2857447|T037|S72.136C|ICD10CM|NONDISPLACED APOPHYSEAL FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP APOPHYSEAL FX UNSP FEMR, INIT FOR OPN FX TYPE 3A/B/C
C2857446|T037|S72.136B|ICD10CM|NONDISPLACED APOPHYSEAL FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP APOPHYSEAL FX UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2848451|T037|S58.919S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED FOREARM, LEVEL UNSPECIFIED, SEQUELA|COMPLETE TRAUMATIC AMP OF UNSP FOREARM, LEVEL UNSP, SEQUELA
C2838223|T037|S32.461B|ICD10CM|DISPLACED ASSOCIATED TRANSVERSE-POSTERIOR FRACTURE OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISPLACED ASSOC TRANSV/POST FX RIGHT ACETAB, INIT FOR OPN FX
C2838222|T037|S32.461A|ICD10CM|DISPLACED ASSOCIATED TRANSVERSE-POSTERIOR FRACTURE OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED ASSOCIATED TRANSV/POST FX RIGHT ACETABULUM, INIT
C2848449|T037|S58.919A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED FOREARM, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMP OF UNSP FOREARM, LEVEL UNSP, INIT
C4237069|T048|F14.980|ICD10CM|COCAINE USE, UNSPECIFIED WITH COCAINE-INDUCED ANXIETY DISORDER|COCAINE INDUCED ANXIETY DISORDER, WITHOUT USE DISORDER
C4237084|T048|F14.981|ICD10CM|COCAINE USE, UNSPECIFIED WITH COCAINE-INDUCED SEXUAL DYSFUNCTION|COCAINE INDUCED SEXUAL DYSFUNCTION, WITHOUT USE DISORDER
C4237087|T048|F14.982|ICD10CM|COCAINE USE, UNSPECIFIED WITH COCAINE-INDUCED SLEEP DISORDER|COCAINE INDUCED SLEEP DISORDER, WITHOUT USE DISORDER
C4268242|T048|F14.988|ICD10CM|COCAINE USE, UNSPECIFIED WITH OTHER COCAINE-INDUCED DISORDER|COCAINE INDUCED OBSESSIVE COMPULSIVE OR RELATED DISORDER
C2887099|T047|A41.89|ICD10CM|OTHER SPECIFIED SEPSIS|OTHER SPECIFIED SEPSIS
C2882217|T047||ICD10CM|SEPTIC PULMONARY EMBOLISM WITH ACUTE COR PULMONALE
C3264366|T047||ICD10CM|SADDLE EMBOLUS OF PULMONARY ARTERY WITH ACUTE COR PULMONALE
C2837766|T037|S32.15XA|ICD10CM|TYPE 2 FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE 2 FRACTURE OF SACRUM, INIT ENCNTR FOR CLOSED FRACTURE
C2882361|T047|I63.29|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF OTHER PRECEREBRAL ARTERIES|CEREBRAL INFRC DUE TO UNSP OCCLS OR STENOSIS OF PRECERB ART
C2837767|T037|S32.15XB|ICD10CM|TYPE 2 FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE 2 FRACTURE OF SACRUM, INIT ENCNTR FOR OPEN FRACTURE
C0588233|T047||ICD10CM|SEPSIS DUE TO ENTEROCOCCUS
C2882218|T047|I26.09|ICD10CM|OTHER PULMONARY EMBOLISM WITH ACUTE COR PULMONALE|OTHER PULMONARY EMBOLISM WITH ACUTE COR PULMONALE
C2902447|T047|M90.569|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, UNSPECIFIED LOWER LEG|OSTEONECROSIS IN DISEASES CLASSD ELSWHR, UNSP LOWER LEG
C2882356|T046|I63.22|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF BASILAR ARTERY|CEREB INFRC DUE TO UNSP OCCLS OR STENOSIS OF BASILAR ARTERY
C2882351|T046|I63.20|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF UNSPECIFIED PRECEREBRAL ARTERIES|CEREB INFRC DUE TO UNSP OCCLS OR STENOS OF UNSP PRECERB ART
C0348642|T047|I68.8|DMDICD10|OTHER CEREBROVASCULAR DISORDERS IN DISEASES CLASSIFIED ELSEWHERE|SONSTIGE ZEREBROVASKULAERE STOERUNGEN BEI ANDERENORTS KLASSIFIZIERTEN KRANKHEITEN
C2921018|T047|E83.118|ICD10CM|OTHER HEMOCHROMATOSIS|OTHER HEMOCHROMATOSIS
C0018995|T047|E83.119|ICD10CM|HEMOCHROMATOSIS, UNSPECIFIED|HEMOCHROMATOSIS, UNSPECIFIED
C0085220|T047|I68.0|DMDICD10|CEREBRAL AMYLOID ANGIOPATHY|ZEREBRALE AMYLOIDANGIOPATHIE
C4290167|T047|I70.55|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF OTHER EXTREMITY WITH ULCERATION|ANY CONDITION CLASSIFIABLE TO I70.518, I70.528, AND I70.538
C2877638|T037|T40.3X2A|ICD10CM|POISONING BY METHADONE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY METHADONE, INTENTIONAL SELF-HARM, INIT ENCNTR
C2921013|T047|E83.110|ICD10CM|HEREDITARY HEMOCHROMATOSIS|PRIMARY (HEREDITARY) HEMOCHROMATOSIS
C2838620|T037|S34.102A|ICD10CM|UNSPECIFIED INJURY TO L2 LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY TO L2 LEVEL OF LUMBAR SPINAL CORD, INIT ENCNTR
C2883736|T037|T50.8X2S|ICD10CM|POISONING BY DIAGNOSTIC AGENTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY DIAGNOSTIC AGENTS, SELF-HARM, SEQUELA
C2877640|T037|T40.3X2S|ICD10CM|POISONING BY METHADONE, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY METHADONE, INTENTIONAL SELF-HARM, SEQUELA
C2856482|T037|S72.001A|ICD10CM|FRACTURE OF UNSPECIFIED PART OF NECK OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF UNSP PART OF NECK OF RIGHT FEMUR, INIT
C2856483|T037|S72.001B|ICD10CM|FRACTURE OF UNSPECIFIED PART OF NECK OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|FX UNSP PART OF NECK OF R FEMUR, INIT FOR OPN FX TYPE I/2
C2856484|T037|S72.001C|ICD10CM|FRACTURE OF UNSPECIFIED PART OF NECK OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|FX UNSP PART OF NECK OF R FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2874524|T048|F13.188|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE WITH OTHER SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED DISORDER|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE W OTH DISORDER
C2874522|T048|F13.181|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED SEXUAL DYSFUNCTION|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE W SEXUAL DYSFUNCTION
C2874521|T048|F13.180|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED ANXIETY DISORDER|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE W ANXIETY DISORDER
C2874523|T048|F13.182|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED SLEEP DISORDER|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE W SLEEP DISORDER
C2882638|T047|I69.865|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING OTHER CEREBROVASCULAR DISEASE, BILATERAL|OTH PARALYTIC SYNDROME FOLLOWING OTH CEREBVASC DISEASE, BI
C2882635|T047|I69.862|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING LEFT DOMINANT SIDE|OTH PARLYT SYND FOL OTH CEREBVASC DISEASE AFF LEFT DOM SIDE
C0752347|T047||ICD10CM|DEMENTIA WITH LEWY BODIES
C4268231|T048|F13.981|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED SEXUAL DYSFUNCTION|SEDATIVE, HYPNOTIC, OR ANXIOLYTIC-INDUCED SEXUAL DYSFUNCTION DISORDER, WITHOUT USE DISORDER
C4237389|T048|F13.232|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH WITHDRAWAL WITH PERCEPTUAL DISTURBANCE|SEDATIVE, HYPNOTIC, OR ANXIOLYTIC WITHDRAWAL WITH PERCEPTUAL DISTURBANCES
C2874535|T048|F13.231|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH WITHDRAWAL DELIRIUM|SEDATV/HYP/ANXIOLYTC DEPENDENCE W WITHDRAWAL DELIRIUM
C2874534|T048|F13.230|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH WITHDRAWAL, UNCOMPLICATED|SEDATV/HYP/ANXIOLYTC DEPENDENCE W WITHDRAWAL, UNCOMPLICATED
C2874175|T047|E13.649|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH HYPOGLYCEMIA WITHOUT COMA|OTH DIABETES MELLITUS WITH HYPOGLYCEMIA WITHOUT COMA
C4237559|T048|F13.988|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH OTHER SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED DISORDER|SEDATIVE, HYPNOTIC, OR ANXIOLYTIC-INDUCED MILD NEUROCOGNITIVE DISORDER
C4237390|T048|F13.239|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE WITH WITHDRAWAL, UNSPECIFIED|SEDATIVE, HYPNOTIC, OR ANXIOLYTIC WITHDRAWAL WITHOUT PERCEPTUAL DISTURBANCES
C0023896|T047|K70|DMDICD10|ALCOHOLIC LIVER DISEASE, UNSPECIFIED|ALKOHOLISCHE LEBERKRANKHEIT
C2874174|T047|E13.641|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH HYPOGLYCEMIA WITH COMA|OTH DIABETES MELLITUS WITH HYPOGLYCEMIA WITH COMA
C2884782|T037|T58.2X2S|ICD10CM|TOXIC EFFECT OF CARBON MONOXIDE FROM INCOMPLETE COMBUSTION OF OTHER DOMESTIC FUELS, INTENTIONAL SELF-HARM, SEQUELA|TOX EFF OF CARB MONX FR INCMPL COMBST DMST FUEL,SLF-HRM,SQLA
C2890821|T037|T84.59XA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO OTHER INTERNAL JOINT PROSTHESIS, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO OTH INTERNAL JOINT PROSTH, INIT
C2835764|T037|S24.103A|ICD10CM|UNSPECIFIED INJURY AT T7-T10 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY AT T7-T10 LEVEL OF THORACIC SPINAL CORD, INIT
C2835765|T037|S24.103D|ICD10CM|UNSPECIFIED INJURY AT T7-T10 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY AT T7-T10 LEVEL OF THORACIC SPINAL CORD, SUBS
C2884780|T037|T58.2X2A|ICD10CM|TOXIC EFFECT OF CARBON MONOXIDE FROM INCOMPLETE COMBUSTION OF OTHER DOMESTIC FUELS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOX EFF OF CARB MONX FR INCMPL COMBST DMST FUEL,SLF-HRM,INIT
C0023944|T047|G83.5|ICD10CM|LOCKED-IN STATE|LOCKED-IN STATE
C4509300|T047|L97.326|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT ANKLE WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULCER OF L ANKLE WITH BONE INVL W/O EVD OF NECR
C4509299|T047|L97.325|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT ANKLE WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULCER OF L ANKLE WITH MSL INVL W/O EVD OF NECR
C2888692|T047|L97.324|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT ANKLE WITH NECROSIS OF BONE|NON-PRESSURE CHRONIC ULCER OF LEFT ANKLE W NECROSIS OF BONE
C2888691|T047|L97.323|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT ANKLE WITH NECROSIS OF MUSCLE|NON-PRS CHRONIC ULCER OF LEFT ANKLE W NECROSIS OF MUSCLE
C2888690|T047|L97.322|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT ANKLE WITH FAT LAYER EXPOSED|NON-PRESSURE CHRONIC ULCER OF LEFT ANKLE W FAT LAYER EXPOSED
C2888689|T047|L97.321|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT ANKLE LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHRONIC ULCER OF LEFT ANKLE LIMITED TO BRKDWN SKIN
C2902729|T047|M96.622|ICD10CM|FRACTURE OF HUMERUS FOLLOWING INSERTION OF ORTHOPEDIC IMPLANT, JOINT PROSTHESIS, OR BONE PLATE, LEFT ARM|FX HUMERUS FOL INSRT ORTHO IMPLNT/PROSTH/BONE PLT, LEFT ARM
C2858869|T037|S72.462B|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL SUPRCNDL FX W INTRCNDL EXTN LOW END L FEMR, 7THB
C2858868|T037|S72.462A|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPL SUPRCNDL FX W INTRCNDL EXTN LOWER END OF L FEMUR, INIT
C0477365|T047|G31.8|ICD10CM|OTHER SPECIFIED DEGENERATIVE DISEASES OF NERVOUS SYSTEM|OTHER SPECIFIED DEGENERATIVE DISEASES OF NERVOUS SYSTEM
C2834056|T037|S14.157A|ICD10CM|OTHER INCOMPLETE LESION AT C7 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|OTH INCOMPLETE LESION AT C7, INIT
C2888693|T047|L97.329|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT ANKLE WITH UNSPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF LEFT ANKLE WITH UNSP SEVERITY
C4509301|T047|L97.328|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT ANKLE WITH OTHER SPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF LEFT ANKLE WITH OTH SEVERITY
C2832515|T037|S06.6X1S|ICD10CM|TRAUMATIC SUBARACHNOID HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|TRAUM SUBRAC HEM W LOC OF 30 MINUTES OR LESS, SEQUELA
C2832399|T037|S06.383A|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF BRAINSTEM WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|CONTUS/LAC/HEM BRAINSTEM W LOC OF 1-5 HRS 59 MIN, INIT
C2883085|T046|I82.221|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF INFERIOR VENA CAVA|CHRONIC EMBOLISM AND THROMBOSIS OF INFERIOR VENA CAVA
C2883084|T046|I82.220|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF INFERIOR VENA CAVA|ACUTE EMBOLISM AND THROMBOSIS OF INFERIOR VENA CAVA
C2901958|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF RIGHT FINGER(S)
C2901959|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF LEFT FINGER(S)
C2901960|T046|M87.046|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED FINGER(S)|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED FINGER(S)
C2901955|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF RIGHT HAND
C2901956|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF LEFT HAND
C2901957|T046|M87.043|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED HAND|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED HAND
C2889352|T047|M05.771|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT ANKLE AND FOOT WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRIT W RHEU FCTR OF RIGHT ANK/FT W/O ORG/SYS INVOLV
C2889353|T047|M05.772|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT ANKLE AND FOOT WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRIT W RHEU FACTOR OF LEFT ANK/FT W/O ORG/SYS INVOLV
C2874378|T048|F10.180|ICD10CM|ALCOHOL ABUSE WITH ALCOHOL-INDUCED ANXIETY DISORDER|ALCOHOL ABUSE WITH ALCOHOL-INDUCED ANXIETY DISORDER
C0268792|T047||ICD10CM|ATHEROEMBOLISM OF KIDNEY
C2874380|T048|F10.182|ICD10CM|ALCOHOL ABUSE WITH ALCOHOL-INDUCED SLEEP DISORDER|ALCOHOL ABUSE WITH ALCOHOL-INDUCED SLEEP DISORDER
C2889354|T047|M05.779|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED ANKLE AND FOOT WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRIT W RHEU FACTOR OF UNSP ANK/FT W/O ORG/SYS INVOLV
C2874381|T048|F10.188|ICD10CM|ALCOHOL ABUSE WITH OTHER ALCOHOL-INDUCED DISORDER|ALCOHOL ABUSE WITH OTHER ALCOHOL-INDUCED DISORDER
C1135216|T047|I75.89|ICD10CM|ATHEROEMBOLISM OF OTHER SITE|ATHEROEMBOLISM OF OTHER SITE
C2833995|T037|S14.141S|ICD10CM|BROWN-SEQUARD SYNDROME AT C1 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|BROWN-SEQUARD SYNDROME AT C1, SEQUELA
C2869880|T037|S98.322S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT MIDFOOT, SEQUELA|PARTIAL TRAUMATIC AMPUTATION OF LEFT MIDFOOT, SEQUELA
C2832545|T037|S06.6X9A|ICD10CM|TRAUMATIC SUBARACHNOID HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|TRAUM SUBRAC HEM W LOC OF UNSP DURATION, INIT
C2837789|T037|S32.19XA|ICD10CM|OTHER FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTHER FRACTURE OF SACRUM, INIT ENCNTR FOR CLOSED FRACTURE
C2869879|T037|S98.322D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT MIDFOOT, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF LEFT MIDFOOT, SUBS ENCNTR
C2833994|T037|S14.141D|ICD10CM|BROWN-SEQUARD SYNDROME AT C1 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|BROWN-SEQUARD SYNDROME AT C1, SUBS
C4268487|T047|I63.433|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF BILATERAL POSTERIOR CEREBRAL ARTERIES|CEREBRAL INFRC DUE TO EMBOLISM OF BI POST CEREBRAL ARTERIES
C2882391|T047|I63.432|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF LEFT POSTERIOR CEREBRAL ARTERY|CEREBRAL INFRC DUE TO EMBOLISM OF LEFT POST CEREBRAL ARTERY
C2882390|T047|I63.431|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF RIGHT POSTERIOR CEREBRAL ARTERY|CEREBRAL INFRC DUE TO EMBOLISM OF RIGHT POST CEREBRAL ARTERY
C2869878|T037|S98.322A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT MIDFOOT, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF LEFT MIDFOOT, INIT ENCNTR
C2832547|T037|S06.6X9S|ICD10CM|TRAUMATIC SUBARACHNOID HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|TRAUM SUBRAC HEM W LOC OF UNSP DURATION, SEQUELA
C2882392|T047|I63.439|ICD10CM|CEREBRAL INFARCTION DUE TO EMBOLISM OF UNSPECIFIED POSTERIOR CEREBRAL ARTERY|CEREBRAL INFRC DUE TO EMBOLISM OF UNSP POST CEREBRAL ARTERY
C2905767|T037|X78.9XXD|ICD10CM|INTENTIONAL SELF-HARM BY UNSPECIFIED SHARP OBJECT, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY UNSP SHARP OBJECT, SUBS ENCNTR
C2837790|T037|S32.19XB|ICD10CM|OTHER FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTHER FRACTURE OF SACRUM, INIT ENCNTR FOR OPEN FRACTURE
C2905766|T037|X78.9XXA|ICD10CM|INTENTIONAL SELF-HARM BY UNSPECIFIED SHARP OBJECT, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY UNSP SHARP OBJECT, INIT ENCNTR
C2859211|T037|S73.031A|ICD10CM|OTHER ANTERIOR SUBLUXATION OF RIGHT HIP, INITIAL ENCOUNTER|OTHER ANTERIOR SUBLUXATION OF RIGHT HIP, INITIAL ENCOUNTER
C4270201|T046|T83.021A|ICD10CM|DISPLACEMENT OF INDWELLING URETHRAL CATHETER, INITIAL ENCOUNTER|DISPLACEMENT OF INDWELLING URETHRAL CATHETER, INIT
C2883308|T037|T49.1X2A|ICD10CM|POISONING BY ANTIPRURITICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ANTIPRURITICS, INTENTIONAL SELF-HARM, INIT
C4236946|T048|F10.988|ICD10CM|ALCOHOL USE, UNSPECIFIED WITH OTHER ALCOHOL-INDUCED DISORDER|ALCOHOL INDUCED MILD NEUROCOGNITIVE DISORDER, WITHOUT USE DISORDER
C2905768|T037|X78.9XXS|ICD10CM|INTENTIONAL SELF-HARM BY UNSPECIFIED SHARP OBJECT, SEQUELA|INTENTIONAL SELF-HARM BY UNSPECIFIED SHARP OBJECT, SEQUELA
C4236934|T048|F10.980|ICD10CM|ALCOHOL USE, UNSPECIFIED WITH ALCOHOL-INDUCED ANXIETY DISORDER|ALCOHOL INDUCED ANXIETY DISORDER, WITHOUT USE DISORDER
C4236952|T048|F10.981|ICD10CM|ALCOHOL USE, UNSPECIFIED WITH ALCOHOL-INDUCED SEXUAL DYSFUNCTION|ALCOHOL INDUCED SEXUAL DYSFUNCTION, WITHOUT USE DISORDER
C4236955|T048|F10.982|ICD10CM|ALCOHOL USE, UNSPECIFIED WITH ALCOHOL-INDUCED SLEEP DISORDER|ALCOHOL INDUCED SLEEP DISORDER, WITHOUT USE DISORDER
C0496763|T191|C08.9|DMDICD10|MALIGNANT NEOPLASM OF MAJOR SALIVARY GLAND, UNSPECIFIED|BOESARTIGE NEUBILDUNG: GROSSE SPEICHELDRUESE, NICHT NAEHER BEZEICHNET
C2890517|T037|T84.053A|ICD10CM|PERIPROSTHETIC OSTEOLYSIS OF INTERNAL PROSTHETIC LEFT KNEE JOINT, INITIAL ENCOUNTER|PERIPROSTH OSTEOLYSIS OF INTERNAL PROSTHETIC L KNEE JT, INIT
C0153361|T191|C08.1|DMDICD10|MALIGNANT NEOPLASM OF SUBLINGUAL GLAND|BOESARTIGE NEUBILDUNG: GLANDULA SUBLINGUALIS
C0153360|T191|C08.0|DMDICD10|MALIGNANT NEOPLASM OF SUBMANDIBULAR GLAND|BOESARTIGE NEUBILDUNG: GLANDULA SUBMANDIBULARIS
C2905804|T037|X82.8XXS|ICD10CM|OTHER INTENTIONAL SELF-HARM BY CRASHING OF MOTOR VEHICLE, SEQUELA|OTH SELF-HARM BY CRASHING OF MOTOR VEHICLE, SEQUELA
C2896619|T046|M80.071A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, RIGHT ANKLE AND FOOT, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, RIGHT ANK/FT, INIT
C2858885|T037|S72.463A|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPL SUPRCNDL FX W INTRCNDL EXTN LOWER END UNSP FEMUR, INIT
C2905803|T037|X82.8XXD|ICD10CM|OTHER INTENTIONAL SELF-HARM BY CRASHING OF MOTOR VEHICLE, SUBSEQUENT ENCOUNTER|OTH INTENTIONAL SELF-HARM BY CRASHING OF MOTOR VEHICLE, SUBS
C2905802|T037|X82.8XXA|ICD10CM|OTHER INTENTIONAL SELF-HARM BY CRASHING OF MOTOR VEHICLE, INITIAL ENCOUNTER|OTH INTENTIONAL SELF-HARM BY CRASHING OF MOTOR VEHICLE, INIT
C4270427|T046|T83.81XA|ICD10CM|EMBOLISM DUE TO GENITOURINARY PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|EMBOLISM DUE TO GENITOURINARY PROSTH DEV/GRFT, INIT
C2838330|T037|S32.484B|ICD10CM|NONDISPLACED DOME FRACTURE OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP DOME FRACTURE OF RIGHT ACETABULUM, INIT FOR OPN FX
C2838329|T037|S32.484A|ICD10CM|NONDISPLACED DOME FRACTURE OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED DOME FRACTURE OF RIGHT ACETABULUM, INIT
C0085677|T047|G62.1|DMDICD10|ALCOHOLIC POLYNEUROPATHY|ALKOHOL-POLYNEUROPATHIE
C0154762|T047|G62.0|DMDICD10|DRUG-INDUCED POLYNEUROPATHY|ARZNEIMITTELINDUZIERTE POLYNEUROPATHIE
C0154763|T047|G62.2|DMDICD10|POLYNEUROPATHY DUE TO OTHER TOXIC AGENTS|POLYNEUROPATHIE DURCH SONSTIGE TOXISCHE AGENZIEN
C2832686|T037|S06.9X3S|ICD10CM|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, SEQUELA|UNSP INTRACRANIAL INJURY W LOC OF 1-5 HRS 59 MIN, SEQUELA
C0442874|T047||ICD10CM|POLYNEUROPATHY, UNSPECIFIED
C2890678|T037|T84.195A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTERNAL FIXATION DEVICE OF LEFT FEMUR, INITIAL ENCOUNTER|MECH COMPL OF INTERNAL FIXATION DEVICE OF LEFT FEMUR, INIT
C2875109|T047|G40.319|ICD10CM|GENERALIZED IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES, INTRACTABLE, WITHOUT STATUS EPILEPTICUS|GENERALIZED IDIOPATHIC EPILEPSY, INTRACTABLE, W/O STAT EPI
C2832684|T037|S06.9X3A|ICD10CM|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|UNSP INTRACRANIAL INJURY W LOC OF 1-5 HRS 59 MIN, INIT
C2875108|T047|G40.311|ICD10CM|GENERALIZED IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES, INTRACTABLE, WITH STATUS EPILEPTICUS|GENERALIZED IDIOPATHIC EPILEPSY, INTRACTABLE, W STAT EPI
C2887454|T047|J45.32|ICD10CM|MILD PERSISTENT ASTHMA WITH STATUS ASTHMATICUS|MILD PERSISTENT ASTHMA WITH STATUS ASTHMATICUS
C2887453|T047||ICD10CM|MILD PERSISTENT ASTHMA WITH (ACUTE) EXACERBATION
C2887452|T047||ICD10CM|MILD PERSISTENT ASTHMA, UNCOMPLICATED
C2884689|T037|T57.3X2A|ICD10CM|TOXIC EFFECT OF HYDROGEN CYANIDE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF HYDROGEN CYANIDE, SELF-HARM, INIT
C2838430|T037|S32.611B|ICD10CM|DISPLACED AVULSION FRACTURE OF RIGHT ISCHIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISPLACED AVULSION FX RIGHT ISCHIUM, INIT FOR OPN FX
C2838429|T037|S32.611A|ICD10CM|DISPLACED AVULSION FRACTURE OF RIGHT ISCHIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED AVULSION FRACTURE OF RIGHT ISCHIUM, INIT
C2860057|T037|S79.002A|ICD10CM|UNSPECIFIED PHYSEAL FRACTURE OF UPPER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP PHYSEAL FRACTURE OF UPPER END OF LEFT FEMUR, INIT
C2977011|T047|I82.5Y9|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF UNSPECIFIED PROXIMAL LOWER EXTREMITY|CHRONIC EMBLSM AND THOMBOS UNSP DEEP VN UNSP PROX LOW EXTRM
C2882993|T047|I70.731|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF THIGH|ATHSCL TYPE OF BYPASS OF THE RIGHT LEG W ULCERATION OF THIGH
C2882994|T047|I70.732|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF CALF|ATHSCL TYPE OF BYPASS OF THE RIGHT LEG W ULCERATION OF CALF
C2882995|T047|I70.733|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF ANKLE|ATHSCL TYPE OF BYPASS OF THE RIGHT LEG W ULCERATION OF ANKLE
C2882997|T047|I70.734|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF HEEL AND MIDFOOT|ATHSCL TYPE OF BYPASS OF RIGHT LEG W ULCER OF HEEL AND MIDFT
C2882999|T047|I70.735|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF OTHER PART OF FOOT|ATHSCL TYPE OF BYPASS OF THE RIGHT LEG W ULCER OTH PRT FOOT
C2883000|T047|I70.738|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF OTHER PART OF LOWER LEG|ATHSCL TYPE OF BYPASS OF RIGHT LEG W ULCER OTH PRT LOW LEG
C2883001|T047|I70.739|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF UNSPECIFIED SITE|ATHSCL TYPE OF BYPASS OF THE RIGHT LEG W ULCER OF UNSP SITE
C2977010|T047|I82.5Y3|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF PROXIMAL LOWER EXTREMITY, BILATERAL|CHR EMBLSM AND THOMBOS UNSP DEEP VEINS OF PROX LOW EXTRM, BI
C2977009|T047|I82.5Y2|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF LEFT PROXIMAL LOWER EXTREMITY|CHR EMBLSM AND THOMBOS UNSP DEEP VN OF LEFT PROX LOW EXTRM
C0261236|T067|E831.0|ICD9CM|DISORDER OF IRON METABOLISM, UNSPECIFIED|BOAT ACC INJ NEC-UNPOWER
C2888914|T047|M00.852|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, LEFT HIP|ARTHRITIS DUE TO OTHER BACTERIA, LEFT HIP
C2845933|T191|C72.31|ICD10CM|MALIGNANT NEOPLASM OF RIGHT OPTIC NERVE|MALIGNANT NEOPLASM OF RIGHT OPTIC NERVE
C2845934|T191|C72.32|ICD10CM|MALIGNANT NEOPLASM OF LEFT OPTIC NERVE|MALIGNANT NEOPLASM OF LEFT OPTIC NERVE
C2888913|T047|M00.851|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, RIGHT HIP|ARTHRITIS DUE TO OTHER BACTERIA, RIGHT HIP
C2856061|T037|S68.624S|ICD10CM|PARTIAL TRAUMATIC TRANSPHALANGEAL AMPUTATION OF RIGHT RING FINGER, SEQUELA|PARTIAL TRAUMATIC TRNSPHAL AMPUTATION OF R RNG FNGR, SEQUELA
C2888915|T047|M00.859|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, UNSPECIFIED HIP|ARTHRITIS DUE TO OTHER BACTERIA, UNSPECIFIED HIP
C2833249|T037|S12.120A|ICD10CM|OTHER DISPLACED DENS FRACTURE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH DISPLACED DENS FRACTURE, INIT ENCNTR FOR CLOSED FRACTURE
C2833250|T037|S12.120B|ICD10CM|OTHER DISPLACED DENS FRACTURE, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTHER DISPLACED DENS FRACTURE, INIT ENCNTR FOR OPEN FRACTURE
C2882315|T047|I60.7|ICD10CM|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM UNSPECIFIED INTRACRANIAL ARTERY|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM UNSP INTRACRAN ART
C2858081|T037|S72.354C|ICD10CM|NONDISPLACED COMMINUTED FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP COMMNT FX SHAFT OF R FEMR, 7THC
C2856518|T037|S72.009C|ICD10CM|FRACTURE OF UNSPECIFIED PART OF NECK OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|FX UNSP PART OF NK OF UNSP FEMR, INIT FOR OPN FX TYPE 3A/B/C
C2858080|T037|S72.354B|ICD10CM|NONDISPLACED COMMINUTED FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP COMMNT FX SHAFT OF R FEMUR, INIT FOR OPN FX TYPE I/2
C2860178|T037|S79.129A|ICD10CM|SALTER-HARRIS TYPE II PHYSEAL FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SLTR-HARIS TYPE II PHYSEAL FX LOWER END OF UNSP FEMUR, INIT
C2858079|T037|S72.354A|ICD10CM|NONDISPLACED COMMINUTED FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP COMMINUTED FRACTURE OF SHAFT OF RIGHT FEMUR, INIT
C2885375|T037|T63.042S|ICD10CM|TOXIC EFFECT OF COBRA VENOM, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF COBRA VENOM, INTENTIONAL SELF-HARM, SEQUELA
C2854074|T191|C88.4|ICD10CM|EXTRANODAL MARGINAL ZONE B-CELL LYMPHOMA OF MUCOSA-ASSOCIATED LYMPHOID TISSUE [MALT-LYMPHOMA]|LYMPHOMA OF SKIN-ASSOCIATED LYMPHOID TISSUE [SALT-LYMPHOMA]
C2854071|T191|C88.0|ICD10CM|WALDENSTROM MACROGLOBULINEMIA|MACROGLOBULINEMIA (IDIOPATHIC) (PRIMARY)
C0021071|T191|C88.3|DMDICD10|IMMUNOPROLIFERATIVE SMALL INTESTINAL DISEASE|IMMUNPROLIFERATIVE DUENNDARMKRANKHEIT
C0242310|T191|C88.2|ICD10CM|HEAVY CHAIN DISEASE|MU HEAVY CHAIN DISEASE
C1264191|T191|C88|DMDICD10|MALIGNANT IMMUNOPROLIFERATIVE DISEASE, UNSPECIFIED|BOESARTIGE IMMUNPROLIFERATIVE KRANKHEITEN
C0348391|T191|C88.8|ICD10CM|OTHER MALIGNANT IMMUNOPROLIFERATIVE DISEASES|OTHER MALIGNANT IMMUNOPROLIFERATIVE DISEASES
C2856088|T037|S68.711S|ICD10CM|COMPLETE TRAUMATIC TRANSMETACARPAL AMPUTATION OF RIGHT HAND, SEQUELA|COMPLETE TRAUMATIC TRANSMETCRPL AMP OF RIGHT HAND, SEQUELA
C2910017|T047|P36.10|ICD10CM|SEPSIS OF NEWBORN DUE TO UNSPECIFIED STREPTOCOCCI|SEPSIS OF NEWBORN DUE TO UNSPECIFIED STREPTOCOCCI
C2888771|T047|L97.929|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF LEFT LOWER LEG WITH UNSPECIFIED SEVERITY|NON-PRS CHRONIC ULC UNSP PRT OF L LOW LEG W UNSP SEVERITY
C4509337|T047|L97.928|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF LEFT LOWER LEG WITH OTHER SPECIFIED SEVERITY|NON-PRS CHRONIC ULC UNSP PRT OF L LOW LEG WITH OTH SEVERITY
C4509335|T047|L97.925|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF LEFT LOWER LEG WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC UNSP PRT L LW LEG W MSL INVL W/O EVD OF NECR
C2888770|T047|L97.924|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF LEFT LOWER LEG WITH NECROSIS OF BONE|NON-PRS CHRONIC ULC UNSP PRT OF L LOW LEG W NECROSIS OF BONE
C4509336|T047|L97.926|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF LEFT LOWER LEG WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC UNSP PRT L LW LEG W BNE INVL W/O EVD OF NECR
C2888767|T047|L97.921|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF LEFT LOWER LEG LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHR ULC UNSP PRT OF L LOW LEG LIMITED TO BRKDWN SKIN
C2888769|T047|L97.923|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF LEFT LOWER LEG WITH NECROSIS OF MUSCLE|NON-PRS CHRONIC ULC UNSP PRT OF L LOW LEG W NECROS MUSCLE
C2888768|T047|L97.922|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF LEFT LOWER LEG WITH FAT LAYER EXPOSED|NON-PRS CHR ULC UNSP PRT OF L LOW LEG W FAT LAYER EXPOSED
C2874825|T048|F19.25|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH PSYCHOACTIVE SUBSTANCE-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH PSYCHOACTIVE SUBSTANCE-INDUCED PSYCHOTIC DISORDER
C2848464|T037|S58.929S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED FOREARM, LEVEL UNSPECIFIED, SEQUELA|PARTIAL TRAUMATIC AMP OF UNSP FOREARM, LEVEL UNSP, SEQUELA
C2890394|T037|T83.89XA|ICD10CM|OTHER SPECIFIED COMPLICATION OF GENITOURINARY PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|OTH COMPLICATION OF GENITOURINARY PROSTH DEV/GRFT, INIT
C2848462|T037|S58.929A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED FOREARM, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP OF UNSP FOREARM, LEVEL UNSP, INIT
C2901930|T047|M86.671|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, RIGHT ANKLE AND FOOT|OTHER CHRONIC OSTEOMYELITIS, RIGHT ANKLE AND FOOT
C2901931|T047|M86.672|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, LEFT ANKLE AND FOOT|OTHER CHRONIC OSTEOMYELITIS, LEFT ANKLE AND FOOT
C2879362|T037|T45.92XA|ICD10CM|POISONING BY UNSPECIFIED PRIMARILY SYSTEMIC AND HEMATOLOGICAL AGENT, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY UNSP PRIM SYS AND HEMATOLOG AGENT, SLF-HRM, INIT
C2901932|T047|M86.679|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, UNSPECIFIED ANKLE AND FOOT|OTHER CHRONIC OSTEOMYELITIS, UNSPECIFIED ANKLE AND FOOT
C2885662|T037|T63.442S|ICD10CM|TOXIC EFFECT OF VENOM OF BEES, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF BEES, SELF-HARM, SEQUELA
C2882360|T046|I63.239|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF UNSPECIFIED CAROTID ARTERIES|CEREB INFRC DUE TO UNSP OCCLS OR STENOS OF UNSP CAROTID ART
C2883111|T047|I82.449|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED TIBIAL VEIN|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED TIBIAL VEIN
C2885660|T037|T63.442A|ICD10CM|TOXIC EFFECT OF VENOM OF BEES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF BEES, INTENTIONAL SELF-HARM, INIT
C2882358|T046|I63.231|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF RIGHT CAROTID ARTERIES|CEREB INFRC DUE TO UNSP OCCLS OR STENOS OF RIGHT CAROTID ART
C2905677|T037|X73.0XXS|ICD10CM|INTENTIONAL SELF-HARM BY SHOTGUN DISCHARGE, SEQUELA|INTENTIONAL SELF-HARM BY SHOTGUN DISCHARGE, SEQUELA
C4268480|T046|I63.233|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF BILATERAL CAROTID ARTERIES|CEREB INFRC DUE TO UNSP OCCLS OR STENOSIS OF BI CAROTID ART
C2882359|T046|I63.232|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF LEFT CAROTID ARTERIES|CEREB INFRC DUE TO UNSP OCCLS OR STENOS OF LEFT CAROTID ART
C2854099|T191||ICD10CM|HAIRY CELL LEUKEMIA NOT HAVING ACHIEVED REMISSION
C0836966|T191||ICD10AM|HAIRY CELL LEUKEMIA, IN REMISSION
C2854100|T191||ICD10CM|HAIRY CELL LEUKEMIA, IN RELAPSE
C4268140|T047|E13.3399|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|OTH DIAB WITH MOD NONP RTNOP WITHOUT MACULAR EDEMA, UNSP
C4268139|T047|E13.3393|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|OTH DIAB WITH MODERATE NONP RTNOP WITHOUT MACULAR EDEMA, BI
C4268138|T047|E13.3392|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|OTH DIAB WITH MOD NONP RTNOP WITHOUT MACULAR EDEMA, L EYE
C4268137|T047|E13.3391|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|OTH DIAB WITH MOD NONP RTNOP WITHOUT MACULAR EDEMA, R EYE
C0837418|T046|M02.19|ICD10CM|POSTDYSENTERIC ARTHROPATHY, MULTIPLE SITES|POSTDYSENTERIC ARTHROPATHY, MULTIPLE SITES
C2889020|T046||ICD10CM|POSTDYSENTERIC ARTHROPATHY, VERTEBRAE
C2832469|T037|S06.5X0A|ICD10CM|TRAUMATIC SUBDURAL HEMORRHAGE WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|TRAUM SUBDR HEM W/O LOSS OF CONSCIOUSNESS, INIT
C0837418|T046|M02.10|ICD10AM|POSTDYSENTERIC ARTHROPATHY, UNSPECIFIED SITE|POSTDYSENTERIC ARTHROPATHY, MULTIPLE SITES
C2832226|T037|S06.341S|ICD10CM|TRAUMATIC HEMORRHAGE OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|TRAUM HEMOR R CEREB W LOC OF 30 MINUTES OR LESS, SEQUELA
C2869772|T037|S98.022A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT FOOT AT ANKLE LEVEL, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP OF LEFT FOOT AT ANKLE LEVEL, INIT
C0282525|T047||ICD10CM|NEONATAL ADRENOLEUKODYSTROPHY
C0043459|T047||ICD10CM|ZELLWEGER SYNDROME
C2832471|T037|S06.5X0S|ICD10CM|TRAUMATIC SUBDURAL HEMORRHAGE WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|TRAUM SUBDR HEM W/O LOSS OF CONSCIOUSNESS, SEQUELA
C2832224|T037|S06.341A|ICD10CM|TRAUMATIC HEMORRHAGE OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|TRAUM HEMOR RIGHT CEREBRUM W LOC OF 30 MINUTES OR LESS, INIT
C2874248|T047|E71.518|ICD10CM|OTHER DISORDERS OF PEROXISOME BIOGENESIS|OTHER DISORDERS OF PEROXISOME BIOGENESIS
C2889987|T037|T82.43XA|ICD10CM|LEAKAGE OF VASCULAR DIALYSIS CATHETER, INITIAL ENCOUNTER|LEAKAGE OF VASCULAR DIALYSIS CATHETER, INITIAL ENCOUNTER
C2833138|T037|S12.000A|ICD10CM|UNSPECIFIED DISPLACED FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP DISP FX OF FIRST CERVICAL VERTEBRA, INIT FOR CLOS FX
C2833139|T037|S12.000B|ICD10CM|UNSPECIFIED DISPLACED FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP DISP FX OF FIRST CERVICAL VERTEBRA, INIT FOR OPN FX
C2855951|T037|S68.412A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT HAND AT WRIST LEVEL, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMP OF LEFT HAND AT WRIST LEVEL, INIT
C2873741|T191||ICD10CM|NEOPLASM OF UNSPECIFIED BEHAVIOR OF BRAIN
C2830286|T047|B66.4|ICD10CM|PARAGONIMIASIS|INFECTION DUE TO PARAGONIMUS SPECIES
C2832674|T037|S06.9X0S|ICD10CM|UNSPECIFIED INTRACRANIAL INJURY WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|UNSP INTRACRANIAL INJURY W/O LOSS OF CONSCIOUSNESS, SEQUELA
C2905668|T037|X71.9XXS|ICD10CM|INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION, UNSPECIFIED, SEQUELA|INTENTIONAL SELF-HARM BY DROWN, UNSP, SEQUELA
C0264323|T047|J42|ICD10CM|UNSPECIFIED CHRONIC BRONCHITIS|CHRONIC TRACHEOBRONCHITIS
C2890787|T037|T84.428A|ICD10CM|DISPLACEMENT OF OTHER INTERNAL ORTHOPEDIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|DISPLACMNT OF INTERNAL ORTH DEVICES, IMPLNT AND GRAFTS, INIT
C2855953|T037|S68.412S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT HAND AT WRIST LEVEL, SEQUELA|COMPLETE TRAUMATIC AMP OF LEFT HAND AT WRIST LEVEL, SEQUELA
C4509310|T047|L97.428|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT HEEL AND MIDFOOT WITH OTHER SPECIFIED SEVERITY|NON-PRS CHRONIC ULCER OF LEFT HEEL/MIDFT WITH OTH SEVERITY
C2833945|T037|S14.127S|ICD10CM|CENTRAL CORD SYNDROME AT C7 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|CENTRAL CORD SYNDROME AT C7, SEQUELA
C2905667|T037|X71.9XXD|ICD10CM|INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION, UNSPECIFIED, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION, UNSP, SUBS
C2832567|T037|S06.814S|ICD10CM|INJURY OF RIGHT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|INJURY OF R INT CAROTID, INTCR W LOC OF 6-24 HRS, SEQUELA
C2837546|T037|S32.029B|ICD10CM|UNSPECIFIED FRACTURE OF SECOND LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF SECOND LUMBAR VERTEBRA, INIT FOR OPN FX
C2888713|T047|L97.429|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT HEEL AND MIDFOOT WITH UNSPECIFIED SEVERITY|NON-PRS CHRONIC ULCER OF LEFT HEEL AND MIDFOOT W UNSP SEVERT
C2832565|T037|S06.814A|ICD10CM|INJURY OF RIGHT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|INJURY OF R INT CAROTID, INTCR W LOC OF 6-24 HRS, INIT
C4269349|T037|S02.32XA|ICD10CM|FRACTURE OF ORBITAL FLOOR, LEFT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF ORBITAL FLOOR, LEFT SIDE, INIT
C2837545|T037|S32.029A|ICD10CM|UNSPECIFIED FRACTURE OF SECOND LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF SECOND LUMBAR VERTEBRA, INIT FOR CLOS FX
C0840027|T037|M87.188|ICD10CM|OSTEONECROSIS DUE TO DRUGS, OTHER SITE|OSTEONECROSIS DUE TO DRUGS, OTHER SITE
C2855968|T037|S68.429A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED HAND AT WRIST LEVEL, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP OF UNSP HAND AT WRIST LEVEL, INIT
C2902031|T047||ICD10CM|OSTEONECROSIS DUE TO DRUGS, JAW
C2833518|T037|S12.500B|ICD10CM|UNSPECIFIED DISPLACED FRACTURE OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP DISP FX OF SIXTH CERVICAL VERTEBRA, INIT FOR OPN FX
C2832431|T037|S06.4X0S|ICD10CM|EPIDURAL HEMORRHAGE WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|EPIDURAL HEMORRHAGE WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA
C2833517|T037|S12.500A|ICD10CM|UNSPECIFIED DISPLACED FRACTURE OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP DISP FX OF SIXTH CERVICAL VERTEBRA, INIT FOR CLOS FX
C2889540|T047|M08.052|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, LEFT HIP|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, LEFT HIP
C2889539|T047|M08.051|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, RIGHT HIP|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, RIGHT HIP
C2889541|T047|M08.059|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED HIP|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED HIP
C2882213|T047|I25.812|ICD10CM|ATHEROSCLEROSIS OF BYPASS GRAFT OF CORONARY ARTERY OF TRANSPLANTED HEART WITHOUT ANGINA PECTORIS|ATHSCL BYPASS OF COR ART OF TRANSPLANTED HEART W/O ANG PCTRS
C2882211|T047|I25.811|ICD10CM|ATHEROSCLEROSIS OF NATIVE CORONARY ARTERY OF TRANSPLANTED HEART WITHOUT ANGINA PECTORIS|ATHSCL NATIVE COR ART OF TRANSPLANTED HEART W/O ANG PCTRS
C2882209|T047|I25.810|ICD10CM|ATHEROSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT(S) WITHOUT ANGINA PECTORIS|ATHEROSCLEROSIS OF CABG W/O ANGINA PECTORIS
C2875321|T047|G72.49|ICD10CM|OTHER INFLAMMATORY AND IMMUNE MYOPATHIES, NOT ELSEWHERE CLASSIFIED|OTH INFLAMMATORY AND IMMUNE MYOPATHIES, NEC
C2869821|T037|S98.141D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF ONE RIGHT LESSER TOE, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF ONE RIGHT LESSER TOE, SUBS
C0238190|T047||ICD10CM|INCLUSION BODY MYOSITIS [IBM]
C2855898|T037|S68.118S|ICD10CM|COMPLETE TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF OTHER FINGER, SEQUELA|COMPLETE TRAUMATIC MCP AMPUTATION OF FINGER, SEQUELA
C2858286|T037|S72.401A|ICD10CM|UNSPECIFIED FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF LOWER END OF RIGHT FEMUR, INIT FOR CLOS FX
C2858287|T037|S72.401B|ICD10CM|UNSPECIFIED FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP FX LOWER END OF RIGHT FEMUR, INIT FOR OPN FX TYPE I/2
C2858288|T037|S72.401C|ICD10CM|UNSPECIFIED FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP FX LOWER END OF R FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2845904|T191|C69.12|ICD10CM|MALIGNANT NEOPLASM OF LEFT CORNEA|MALIGNANT NEOPLASM OF LEFT CORNEA
C2837954|T191|C34.30|ICD10CM|MALIGNANT NEOPLASM OF LOWER LOBE, UNSPECIFIED BRONCHUS OR LUNG|MALIGNANT NEOPLASM OF LOWER LOBE, UNSP BRONCHUS OR LUNG
C2845903|T191|C69.11|ICD10CM|MALIGNANT NEOPLASM OF RIGHT CORNEA|MALIGNANT NEOPLASM OF RIGHT CORNEA
C2889108|T047|M05.011|ICD10CM|FELTY'S SYNDROME, RIGHT SHOULDER|FELTY'S SYNDROME, RIGHT SHOULDER
C2889109|T047|M05.012|ICD10CM|FELTY'S SYNDROME, LEFT SHOULDER|FELTY'S SYNDROME, LEFT SHOULDER
C2889110|T047|M05.019|ICD10CM|FELTY'S SYNDROME, UNSPECIFIED SHOULDER|FELTY'S SYNDROME, UNSPECIFIED SHOULDER
C2888949|T047|M01.X59|ICD10CM|DIRECT INFECTION OF UNSPECIFIED HIP IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIRECT INFCT OF UNSP HIP IN INFEC/PARASTC DIS CLASSD ELSWHR
C2835233|T037|S22.021A|ICD10CM|STABLE BURST FRACTURE OF SECOND THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|STABLE BURST FRACTURE OF SECOND THORACIC VERTEBRA, INIT
C2835234|T037|S22.021B|ICD10CM|STABLE BURST FRACTURE OF SECOND THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|STABLE BURST FX SECOND THOR VERTEBRA, INIT FOR OPN FX
C2888947|T047|M01.X51|ICD10CM|DIRECT INFECTION OF RIGHT HIP IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIRECT INFCT OF R HIP IN INFEC/PARASTC DIS CLASSD ELSWHR
C2837517|T037|S32.020A|ICD10CM|WEDGE COMPRESSION FRACTURE OF SECOND LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|WEDGE COMPRESSION FRACTURE OF SECOND LUMBAR VERTEBRA, INIT
C2888948|T047|M01.X52|ICD10CM|DIRECT INFECTION OF LEFT HIP IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIRECT INFCT OF LEFT HIP IN INFEC/PARASTC DIS CLASSD ELSWHR
C4269434|T037|S02.602B|ICD10CM|FRACTURE OF UNSPECIFIED PART OF BODY OF LEFT MANDIBLE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF UNSPECIFIED PART OF BODY OF LEFT MANDIBLE, 7THB
C2869822|T037|S98.141S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF ONE RIGHT LESSER TOE, SEQUELA|PARTIAL TRAUMATIC AMP OF ONE RIGHT LESSER TOE, SEQUELA
C4269433|T037|S02.602A|ICD10CM|FRACTURE OF UNSPECIFIED PART OF BODY OF LEFT MANDIBLE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF UNSPECIFIED PART OF BODY OF LEFT MANDIBLE, INIT
C2885390|T037|T63.062A|ICD10CM|TOXIC EFFECT OF VENOM OF OTHER NORTH AND SOUTH AMERICAN SNAKE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF N & S AMERICAN SNAKE, SLF-HRM, INIT
C2857701|T037|S72.309A|ICD10CM|UNSPECIFIED FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF SHAFT OF UNSP FEMUR, INIT FOR CLOS FX
C2857703|T037|S72.309C|ICD10CM|UNSPECIFIED FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP FX SHAFT OF UNSP FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2857702|T037|S72.309B|ICD10CM|UNSPECIFIED FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP FX SHAFT OF UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2837684|T037|S32.112B|ICD10CM|SEVERELY DISPLACED ZONE I FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|SEVERELY DISPLACED ZONE I FX SACRUM, INIT FOR OPN FX
C2837683|T037|S32.112A|ICD10CM|SEVERELY DISPLACED ZONE I FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SEVERELY DISPLACED ZONE I FRACTURE OF SACRUM, INIT
C4269438|T037|S02.602S|ICD10CM|FRACTURE OF UNSPECIFIED PART OF BODY OF LEFT MANDIBLE, SEQUELA|FX UNSPECIFIED PART OF BODY OF LEFT MANDIBLE, SEQUELA
C2885392|T037|T63.062S|ICD10CM|TOXIC EFFECT OF VENOM OF OTHER NORTH AND SOUTH AMERICAN SNAKE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF N & S AMERICAN SNAKE, SLF-HRM, SQLA
C2879723|T037|T47.2X2S|ICD10CM|POISONING BY STIMULANT LAXATIVES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY STIMULANT LAXATIVES, SELF-HARM, SEQUELA
C0264332|T046||ICD10CM|TRACHEO-ESOPHAGEAL FISTULA FOLLOWING TRACHEOSTOMY
C2838637|T037|S34.109D|ICD10CM|UNSPECIFIED INJURY TO UNSPECIFIED LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY TO UNSP LEVEL OF LUMBAR SPINAL CORD, SUBS ENCNTR
C2838636|T037|S34.109A|ICD10CM|UNSPECIFIED INJURY TO UNSPECIFIED LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY TO UNSP LEVEL OF LUMBAR SPINAL CORD, INIT ENCNTR
C4270552|T046|T85.635A|ICD10CM|LEAKAGE OF OTHER NERVOUS SYSTEM DEVICE, IMPLANT OR GRAFT, INITIAL ENCOUNTER|LEAKAGE OF OTHER NERVOUS SYS DEVICE, IMPLANT OR GRAFT, INIT
C2879721|T037|T47.2X2A|ICD10CM|POISONING BY STIMULANT LAXATIVES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY STIMULANT LAXATIVES, SELF-HARM, INIT
C2832610|T037|S06.825A|ICD10CM|INJURY OF LEFT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, INITIAL ENCOUNTER|INJ L INT CAROTID, INTCR W LOC >24 HR W RET CONSC LEV, INIT
C2838638|T037|S34.109S|ICD10CM|UNSPECIFIED INJURY TO UNSPECIFIED LEVEL OF LUMBAR SPINAL CORD, SEQUELA|UNSP INJURY TO UNSP LEVEL OF LUMBAR SPINAL CORD, SEQUELA
C2886347|T037|T71.122A|ICD10CM|ASPHYXIATION DUE TO PLASTIC BAG, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|ASPHYXIATION DUE TO PLASTIC BAG, INTENTIONAL SELF-HARM, INIT
C0349049|T191|C16.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF STOMACH|BOESARTIGE NEUBILDUNG: MAGEN, MEHRERE TEILBEREICHE UEBERLAPPEND
C0024623|T191|C16.9|DMDICD10|MALIGNANT NEOPLASM OF STOMACH, UNSPECIFIED|BOESARTIGE NEUBILDUNG: MAGEN, NICHT NAEHER BEZEICHNET
C2837935|T191|C16.6|ICD10CM|MALIGNANT NEOPLASM OF GREATER CURVATURE OF STOMACH, UNSPECIFIED|MALIGNANT NEOPLASM OF GREATER CURVATURE OF STOMACH, NOT CLASSIFIABLE TO C16.0-C16.4
C0153418|T191|C16.4|DMDICD10|MALIGNANT NEOPLASM OF PYLORUS|BOESARTIGE NEUBILDUNG: PYLORUS
C2837934|T191|C16.5|ICD10CM|MALIGNANT NEOPLASM OF LESSER CURVATURE OF STOMACH, UNSPECIFIED|MALIGNANT NEOPLASM OF LESSER CURVATURE OF STOMACH, NOT CLASSIFIABLE TO C16.1-C16.4
C0153421|T191|C16.2|DMDICD10|MALIGNANT NEOPLASM OF BODY OF STOMACH|BOESARTIGE NEUBILDUNG: CORPUS VENTRICULI
C2837933|T191|C16.3|ICD10CM|MALIGNANT NEOPLASM OF PYLORIC ANTRUM|MALIGNANT NEOPLASM OF GASTRIC ANTRUM
C2837932|T191|C16.0|ICD10CM|MALIGNANT NEOPLASM OF CARDIA|MALIGNANT NEOPLASM OF ESOPHAGUS AND STOMACH
C0153420|T191|C16.1|DMDICD10|MALIGNANT NEOPLASM OF FUNDUS OF STOMACH|BOESARTIGE NEUBILDUNG: FUNDUS VENTRICULI
C2902044|T046|M87.233|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA OF UNSPECIFIED RADIUS|OSTEONECROSIS DUE TO PREVIOUS TRAUMA OF UNSPECIFIED RADIUS
C2902043|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA OF LEFT RADIUS
C2902042|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA OF RIGHT RADIUS
C2902048|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA OF RIGHT CARPUS
C2902047|T046|M87.236|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA OF UNSPECIFIED ULNA|OSTEONECROSIS DUE TO PREVIOUS TRAUMA OF UNSPECIFIED ULNA
C2902046|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA OF LEFT ULNA
C2902045|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA OF RIGHT ULNA
C2902050|T046|M87.239|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA OF UNSPECIFIED CARPUS|OSTEONECROSIS DUE TO PREVIOUS TRAUMA OF UNSPECIFIED CARPUS
C2902049|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA OF LEFT CARPUS
C2856794|T037|S72.041B|ICD10CM|DISPLACED FRACTURE OF BASE OF NECK OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF BASE OF NECK OF R FEMUR, INIT FOR OPN FX TYPE I/2
C2885123|T037|T61.02XA|ICD10CM|CIGUATERA FISH POISONING, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|CIGUATERA FISH POISONING, INTENTIONAL SELF-HARM, INIT ENCNTR
C2875085|T047|G40.109|ICD10CM|LOCALIZATION-RELATED (FOCAL) (PARTIAL) SYMPTOMATIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SIMPLE PARTIAL SEIZURES, NOT INTRACTABLE, WITHOUT STATUS EPILEPTICUS|LOCAL-REL SYMPTC EPI W SIMP PRT SEIZ,NOT NTRCT, W/O STAT EPI
C2838164|T037|S32.445A|ICD10CM|NONDISPLACED FRACTURE OF POSTERIOR COLUMN [ILIOISCHIAL] OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF POSTERIOR COLUMN OF LEFT ACETABULUM, INIT
C2838165|T037|S32.445B|ICD10CM|NONDISPLACED FRACTURE OF POSTERIOR COLUMN [ILIOISCHIAL] OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP FX OF POST COLUMN OF LEFT ACETAB, INIT FOR OPN FX
C2875084|T047|G40.101|ICD10CM|LOCALIZATION-RELATED (FOCAL) (PARTIAL) SYMPTOMATIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SIMPLE PARTIAL SEIZURES, NOT INTRACTABLE, WITH STATUS EPILEPTICUS|LOCAL-REL SYMPTC EPI W SIMP PART SEIZ, NOT NTRCT, W STAT EPI
C2885125|T037|T61.02XS|ICD10CM|CIGUATERA FISH POISONING, INTENTIONAL SELF-HARM, SEQUELA|CIGUATERA FISH POISONING, INTENTIONAL SELF-HARM, SEQUELA
C2902893|T047|N04.8|ICD10CM|NEPHROTIC SYNDROME WITH OTHER MORPHOLOGIC CHANGES|NEPHROTIC SYNDROME WITH OTHER MORPHOLOGIC CHANGES
C2902894|T047|N04.9|ICD10CM|NEPHROTIC SYNDROME WITH UNSPECIFIED MORPHOLOGIC CHANGES|NEPHROTIC SYNDROME WITH UNSPECIFIED MORPHOLOGIC CHANGES
C0451721|T047|N04.2|DMDICD10|NEPHROTIC SYNDROME WITH DIFFUSE MEMBRANOUS GLOMERULONEPHRITIS|NEPHROTISCHES SYNDROM: DIFFUSE MEMBRANOESE GLOMERULONEPHRITIS
C0451722|T047|N04.3|DMDICD10|NEPHROTIC SYNDROME WITH DIFFUSE MESANGIAL PROLIFERATIVE GLOMERULONEPHRITIS|NEPHROTISCHES SYNDROM: DIFFUSE MESANGIOPROLIFERATIVE GLOMERULONEPHRITIS
C2902886|T047|N04.0|ICD10CM|NEPHROTIC SYNDROME WITH MINOR GLOMERULAR ABNORMALITY|NEPHROTIC SYNDROME WITH MINIMAL CHANGE LESION
C2902889|T047|N04.1|ICD10CM|NEPHROTIC SYNDROME WITH FOCAL AND SEGMENTAL GLOMERULAR LESIONS|NEPHROTIC SYNDROME WITH FOCAL GLOMERULONEPHRITIS
C2902891|T047|N04.6|ICD10CM|NEPHROTIC SYNDROME WITH DENSE DEPOSIT DISEASE|NEPHROTIC SYNDROME WITH MEMBRANOPROLIFERATIVE GLOMERULONEPHRITIS, TYPE 2
C2902892|T047|N04.7|ICD10CM|NEPHROTIC SYNDROME WITH DIFFUSE CRESCENTIC GLOMERULONEPHRITIS|NEPHROTIC SYNDROME WITH EXTRACAPILLARY GLOMERULONEPHRITIS
C0451723|T047|N04.4|DMDICD10|NEPHROTIC SYNDROME WITH DIFFUSE ENDOCAPILLARY PROLIFERATIVE GLOMERULONEPHRITIS|NEPHROTISCHES SYNDROM: DIFFUSE ENDOKAPILLAER-PROLIFERATIVE GLOMERULONEPHRITIS
C2902890|T047|N04.5|ICD10CM|NEPHROTIC SYNDROME WITH DIFFUSE MESANGIOCAPILLARY GLOMERULONEPHRITIS|NEPHROTIC SYNDROME WITH MEMBRANOPROLIFERATIVE GLOMERULONEPHRITIS, TYPES 1 AND 3, OR NOS
C2884659|T037|T57.1X2S|ICD10CM|TOXIC EFFECT OF PHOSPHORUS AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF PHOSPHORUS AND ITS COMPND, SLF-HRM, SEQUELA
C2884643|T037|T57.0X2S|ICD10CM|TOXIC EFFECT OF ARSENIC AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF ARSENIC AND ITS COMPND, SELF-HARM, SEQUELA
C2886085|T037|T65.4X2A|ICD10CM|TOXIC EFFECT OF CARBON DISULFIDE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CARBON DISULFIDE, SELF-HARM, INIT
C2884657|T037|T57.1X2A|ICD10CM|TOXIC EFFECT OF PHOSPHORUS AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF PHOSPHORUS AND ITS COMPND, SELF-HARM, INIT
C2884641|T037|T57.0X2A|ICD10CM|TOXIC EFFECT OF ARSENIC AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF ARSENIC AND ITS COMPOUNDS, SELF-HARM, INIT
C2856036|T037|S68.618S|ICD10CM|COMPLETE TRAUMATIC TRANSPHALANGEAL AMPUTATION OF OTHER FINGER, SEQUELA|COMPLETE TRAUMATIC TRNSPHAL AMPUTATION OF FINGER, SEQUELA
C1398892|T047||ICD10CM|GONOCOCCAL SEPSIS
C0018077|T047|A54.85|ICD10CM|GONOCOCCAL PERITONITIS|GONOCOCCAL PERITONITIS
C2893395|T047|A54.84|ICD10CM|GONOCOCCAL PNEUMONIA|GONOCOCCAL PNEUMONIA
C1404114|T046|T86.32|ICD10CM|HEART-LUNG TRANSPLANT FAILURE|HEART-LUNG TRANSPLANT FAILURE
C2891278|T046|T86.33|ICD10CM|HEART-LUNG TRANSPLANT INFECTION|HEART-LUNG TRANSPLANT INFECTION
C2891277|T037|T86.30|ICD10CM|UNSPECIFIED COMPLICATION OF HEART-LUNG TRANSPLANT|UNSPECIFIED COMPLICATION OF HEART-LUNG TRANSPLANT
C0854432|T046|T86.31|ICD10CM|HEART-LUNG TRANSPLANT REJECTION|HEART-LUNG TRANSPLANT REJECTION
C2869908|T037|S98.929A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED FOOT, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF UNSP FOOT, LEVEL UNSP, INIT
C2901321|T046|M84.572A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, LEFT ANKLE, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, LEFT ANKLE, INIT
C2891279|T037|T86.39|ICD10CM|OTHER COMPLICATIONS OF HEART-LUNG TRANSPLANT|OTHER COMPLICATIONS OF HEART-LUNG TRANSPLANT
C2869909|T037|S98.929D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED FOOT, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF UNSP FOOT, LEVEL UNSP, SUBS
C2874295|T047|E80.21|ICD10CM|ACUTE INTERMITTENT (HEPATIC) PORPHYRIA|ACUTE INTERMITTENT (HEPATIC) PORPHYRIA
C2843338|T037|S48.922A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT SHOULDER AND UPPER ARM, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP OF LEFT SHLDR/UP ARM, LEVEL UNSP, INIT
C2857909|T037|S72.336C|ICD10CM|NONDISPLACED OBLIQUE FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP OBLIQUE FX SHAFT OF UNSP FEMR, 7THC
C2869910|T037|S98.929S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED FOOT, LEVEL UNSPECIFIED, SEQUELA|PARTIAL TRAUMATIC AMP OF UNSP FOOT, LEVEL UNSP, SEQUELA
C4270375|T046|T83.712A|ICD10CM|EROSION OF IMPLANTED URETHRAL MESH TO SURROUNDING ORGAN OR TISSUE, INITIAL ENCOUNTER|EROSN IMPLNT URETHRAL MESH TO SURRND ORG/TISS, INIT
C2857908|T037|S72.336B|ICD10CM|NONDISPLACED OBLIQUE FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP OBLIQUE FX SHAFT OF UNSP FEMR, 7THB
C0477468|T047|L10.8|ICD10CM|OTHER PEMPHIGUS|OTHER PEMPHIGUS
C2857907|T037|S72.336A|ICD10CM|NONDISPLACED OBLIQUE FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED OBLIQUE FRACTURE OF SHAFT OF UNSP FEMUR, INIT
C2869811|T037|S98.132A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF ONE LEFT LESSER TOE, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF ONE LEFT LESSER TOE, INIT
C4269326|T037|S02.11GS|ICD10CM|OTHER FRACTURE OF OCCIPUT, RIGHT SIDE, SEQUELA|OTHER FRACTURE OF OCCIPUT, RIGHT SIDE, SEQUELA
C1112570|T191|L10.81|ICD10CM|PARANEOPLASTIC PEMPHIGUS|PARANEOPLASTIC PEMPHIGUS
C2869812|T037|S98.132D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF ONE LEFT LESSER TOE, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF ONE LEFT LESSER TOE, SUBS
C4269321|T037|S02.11GA|ICD10CM|OTHER FRACTURE OF OCCIPUT, RIGHT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTHER FRACTURE OF OCCIPUT, RIGHT SIDE, INIT
C2869813|T037|S98.132S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF ONE LEFT LESSER TOE, SEQUELA|COMPLETE TRAUMATIC AMP OF ONE LEFT LESSER TOE, SEQUELA
C4269322|T037|S02.11GB|ICD10CM|OTHER FRACTURE OF OCCIPUT, RIGHT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTHER FRACTURE OF OCCIPUT, RIGHT SIDE, 7THB
C2874980|T048|F63.9|ICD10CM|IMPULSE DISORDER, UNSPECIFIED|IMPULSE DISORDER, UNSPECIFIED
C0348496|T047|E80.29|ICD10CM|OTHER PORPHYRIA|OTHER PORPHYRIA
C0016142|T048|F63.1|DMDICD10|PYROMANIA|PATHOLOGISCHE BRANDSTIFTUNG [PYROMANIE]
C0030662|T048|F63.0|DMDICD10|PATHOLOGICAL GAMBLING|PATHOLOGISCHES SPIELEN
C0040953|T048|F63.3|DMDICD10|TRICHOTILLOMANIA|TRICHOTILLOMANIE
C0022734|T048|F63.2|DMDICD10|KLEPTOMANIA|PATHOLOGISCHES STEHLEN [KLEPTOMANIE]
C2833219|T037|S12.101A|ICD10CM|UNSPECIFIED NONDISPLACED FRACTURE OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP NONDISP FX OF SECOND CERVICAL VERTEBRA, INIT
C2833220|T037|S12.101B|ICD10CM|UNSPECIFIED NONDISPLACED FRACTURE OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP NONDISP FX OF SECOND CERVICAL VERTEBRA, INIT FOR OPN FX
C2879053|T037|T45.1X2S|ICD10CM|POISONING BY ANTINEOPLASTIC AND IMMUNOSUPPRESSIVE DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY ANTINEOPL AND IMMUNOSUP DRUGS, SELF-HARM, SEQUELA
C2884272|T037|T53.4X2S|ICD10CM|TOXIC EFFECT OF DICHLOROMETHANE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF DICHLOROMETHANE, SELF-HARM, SEQUELA
C2838336|T037|S32.485A|ICD10CM|NONDISPLACED DOME FRACTURE OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED DOME FRACTURE OF LEFT ACETABULUM, INIT
C2879026|T037|T45.0X2A|ICD10CM|POISONING BY ANTIALLERGIC AND ANTIEMETIC DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ANTIALLERG/ANTIEMETIC, SELF-HARM, INIT
C2886457|T037|T71.222A|ICD10CM|ASPHYXIATION DUE TO BEING TRAPPED IN A CAR TRUNK, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|ASPHYX DUE TO BEING TRAPPED IN A CAR TRUNK, SELF-HARM, INIT
C2838337|T037|S32.485B|ICD10CM|NONDISPLACED DOME FRACTURE OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP DOME FRACTURE OF LEFT ACETABULUM, INIT FOR OPN FX
C2911488|T033|Z93.50|ICD10CM|UNSPECIFIED CYSTOSTOMY STATUS|UNSPECIFIED CYSTOSTOMY STATUS
C2911489|T033|Z93.51|ICD10CM|CUTANEOUS-VESICOSTOMY STATUS|CUTANEOUS-VESICOSTOMY STATUS
C2879051|T037|T45.1X2A|ICD10CM|POISONING BY ANTINEOPLASTIC AND IMMUNOSUPPRESSIVE DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ANTINEOPL AND IMMUNOSUP DRUGS, SELF-HARM, INIT
C2884270|T037|T53.4X2A|ICD10CM|TOXIC EFFECT OF DICHLOROMETHANE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF DICHLOROMETHANE, INTENTIONAL SELF-HARM, INIT
C2896713|T046|M80.832A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, LEFT FOREARM, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, L FOREARM, INIT
C0040517|T047|F95.2|DMDICD10|TOURETTE'S DISORDER|KOMBINIERTE VOKALE UND MULTIPLE MOTORISCHE TICS [TOURETTE-SYNDROM]
C2911491|T033|Z93.59|ICD10CM|OTHER CYSTOSTOMY STATUS|OTHER CYSTOSTOMY STATUS
C2879028|T037|T45.0X2S|ICD10CM|POISONING BY ANTIALLERGIC AND ANTIEMETIC DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ANTIALLERG/ANTIEMETIC, SELF-HARM, SEQUELA
C2886459|T037|T71.222S|ICD10CM|ASPHYXIATION DUE TO BEING TRAPPED IN A CAR TRUNK, INTENTIONAL SELF-HARM, SEQUELA|ASPHYX DUE TO BEING TRAPPED IN A CAR TRUNK, SLF-HRM, SEQUELA
C3250150|T047|E05.41|ICD10CM|THYROTOXICOSIS FACTITIA WITH THYROTOXIC CRISIS OR STORM|THYROTOXICOSIS FACTITIA WITH THYROTOXIC CRISIS OR STORM
C2873873|T047||ICD10CM|THYROTOXICOSIS FACTITIA WITHOUT THYROTOXIC CRISIS OR STORM
C2889478|T047|M06.841|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, RIGHT HAND|OTHER SPECIFIED RHEUMATOID ARTHRITIS, RIGHT HAND
C2889480|T047|M06.849|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, UNSPECIFIED HAND|OTHER SPECIFIED RHEUMATOID ARTHRITIS, UNSPECIFIED HAND
C2362742|T019|Q04.3|ICD10CM|OTHER REDUCTION DEFORMITIES OF BRAIN|MICROGYRIA
C0079541|T019|Q04.2|DMDICD10|HOLOPROSENCEPHALY|HOLOPROSENZEPHALIE-SYNDROM
C0078982|T019|Q04.1|DMDICD10|ARHINENCEPHALY|ARRHINENZEPHALIE
C0431366|T019|Q04.0|DMDICD10|CONGENITAL MALFORMATIONS OF CORPUS CALLOSUM|ANGEBORENE FEHLBILDUNGEN DES CORPUS CALLOSUM
C0302892|T019|Q04.6|ICD10CM|CONGENITAL CEREBRAL CYSTS|PORENCEPHALY
C2720434|T019|Q04.5|DMDICD10|MEGALENCEPHALY|MEGALENZEPHALIE
C2910099|T019|Q04.4|ICD10CM|SEPTO-OPTIC DYSPLASIA OF BRAIN|SEPTO-OPTIC DYSPLASIA OF BRAIN
C2910102|T019|Q04.9|ICD10CM|CONGENITAL MALFORMATION OF BRAIN, UNSPECIFIED|MULTIPLE ANOMALIES NOS OF BRAIN, CONGENITAL
C2910100|T047|Q04.8|ICD10CM|OTHER SPECIFIED CONGENITAL MALFORMATIONS OF BRAIN|ARNOLD-CHIARI SYNDROME, TYPE IV
C2890834|T037|T84.611A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL FIXATION DEVICE OF LEFT HUMERUS, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INT FIX OF LEFT HUMERUS, INIT
C2977068|T047|J96.11|ICD10CM|CHRONIC RESPIRATORY FAILURE WITH HYPOXIA|CHRONIC RESPIRATORY FAILURE WITH HYPOXIA
C2977067|T047|J96.10|ICD10CM|CHRONIC RESPIRATORY FAILURE, UNSPECIFIED WHETHER WITH HYPOXIA OR HYPERCAPNIA|CHRONIC RESPIRATORY FAILURE, UNSP W HYPOXIA OR HYPERCAPNIA
C2977069|T047|J96.12|ICD10CM|CHRONIC RESPIRATORY FAILURE WITH HYPERCAPNIA|CHRONIC RESPIRATORY FAILURE WITH HYPERCAPNIA
C2856913|T037|S72.052A|ICD10CM|UNSPECIFIED FRACTURE OF HEAD OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF HEAD OF LEFT FEMUR, INIT FOR CLOS FX
C2856914|T037|S72.052B|ICD10CM|UNSPECIFIED FRACTURE OF HEAD OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP FX HEAD OF LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C2856915|T037|S72.052C|ICD10CM|UNSPECIFIED FRACTURE OF HEAD OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP FX HEAD OF LEFT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C4269238|T037|S02.102B|ICD10CM|FRACTURE OF BASE OF SKULL, LEFT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF BASE OF SKULL, LEFT SIDE, 7THB
C4269237|T037|S02.102A|ICD10CM|FRACTURE OF BASE OF SKULL, LEFT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF BASE OF SKULL, LEFT SIDE, INIT
C2842140|T191|C50.921|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF RIGHT MALE BREAST|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF RIGHT MALE BREAST
C2842141|T191|C50.922|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF LEFT MALE BREAST|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF LEFT MALE BREAST
C2875185|T047|G43.901|ICD10CM|MIGRAINE, UNSPECIFIED, NOT INTRACTABLE, WITH STATUS MIGRAINOSUS|MIGRAINE, UNSP, NOT INTRACTABLE, WITH STATUS MIGRAINOSUS
C0475531|T046|D64.2|DMDICD10|SECONDARY SIDEROBLASTIC ANEMIA DUE TO DRUGS AND TOXINS|SEKUNDAERE SIDEROACHRESTISCHE [SIDEROBLASTISCHE] ANAEMIE DURCH ARZNEIMITTEL ODER TOXINE
C2873781|T047|D64.3|ICD10CM|OTHER SIDEROBLASTIC ANEMIAS|PYRIDOXINE-RESPONSIVE SIDEROBLASTIC ANEMIA NEC
C0221018|T047|D64.0|DMDICD10|HEREDITARY SIDEROBLASTIC ANEMIA|HEREDITAERE SIDEROACHRESTISCHE [SIDEROBLASTISCHE] ANAEMIE
C0475532|T047|D64.1|DMDICD10|SECONDARY SIDEROBLASTIC ANEMIA DUE TO DISEASE|SEKUNDAERE SIDEROACHRESTISCHE [SIDEROBLASTISCHE] ANAEMIE (KRANKHEITSBEDINGT)
C4269242|T037|S02.102S|ICD10CM|FRACTURE OF BASE OF SKULL, LEFT SIDE, SEQUELA|FRACTURE OF BASE OF SKULL, LEFT SIDE, SEQUELA
C2875186|T047|G43.909|ICD10CM|MIGRAINE, UNSPECIFIED, NOT INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|MIGRAINE, UNSP, NOT INTRACTABLE, WITHOUT STATUS MIGRAINOSUS
C2857583|T037|S72.22XC|ICD10CM|DISPLACED SUBTROCHANTERIC FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPLACED SUBTROCHNT FX L FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2901794|T047|M86.111|ICD10CM|OTHER ACUTE OSTEOMYELITIS, RIGHT SHOULDER|OTHER ACUTE OSTEOMYELITIS, RIGHT SHOULDER
C0837617|T047|M06.80|ICD10AM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, UNSPECIFIED SITE|OTHER SPECIFIED RHEUMATOID ARTHRITIS, MULTIPLE SITES
C2901795|T047|M86.112|ICD10CM|OTHER ACUTE OSTEOMYELITIS, LEFT SHOULDER|OTHER ACUTE OSTEOMYELITIS, LEFT SHOULDER
C2843314|T037|S48.122S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN LEFT SHOULDER AND ELBOW, SEQUELA|PARTIAL TRAUM AMP AT LEVEL BETW L SHLDR AND ELBOW, SEQUELA
C2901796|T047|M86.119|ICD10CM|OTHER ACUTE OSTEOMYELITIS, UNSPECIFIED SHOULDER|OTHER ACUTE OSTEOMYELITIS, UNSPECIFIED SHOULDER
C2889492|T047|M06.88|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, VERTEBRAE|OTHER SPECIFIED RHEUMATOID ARTHRITIS, VERTEBRAE
C0837617|T047|M06.89|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, MULTIPLE SITES|OTHER SPECIFIED RHEUMATOID ARTHRITIS, MULTIPLE SITES
C2874170|T047|E13.628|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH OTHER SKIN COMPLICATIONS|OTH DIABETES MELLITUS WITH OTHER SKIN COMPLICATIONS
C2874168|T047|E13.621|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH FOOT ULCER|OTHER SPECIFIED DIABETES MELLITUS WITH FOOT ULCER
C2874167|T047|E13.620|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC DERMATITIS|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC DERMATITIS
C2874169|T047|E13.622|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH OTHER SKIN ULCER|OTHER SPECIFIED DIABETES MELLITUS WITH OTHER SKIN ULCER
C0020541|T047|K76.6|DMDICD10|PORTAL HYPERTENSION|PORTALE HYPERTONIE
C0019212|T047|K76.7|DMDICD10|HEPATORENAL SYNDROME|HEPATORENALES SYNDROM
C4290177|T047|I70.75|ICD10CM|ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF OTHER EXTREMITY WITH ULCERATION|ANY CONDITION CLASSIFIABLE TO I70.718 AND I70.728
C2889294|T047|M05.579|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP ANK/FT
C2835854|T037|S24.154D|ICD10CM|OTHER INCOMPLETE LESION AT T11-T12 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|OTH INCOMPLETE LESION AT T11-T12, SUBS
C2835756|T037|S24.101A|ICD10CM|UNSPECIFIED INJURY AT T1 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY AT T1 LEVEL OF THORACIC SPINAL CORD, INIT ENCNTR
C2889293|T047|M05.572|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF LEFT ANK/FT
C2835853|T037|S24.154A|ICD10CM|OTHER INCOMPLETE LESION AT T11-T12 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|OTH INCOMPLETE LESION AT T11-T12, INIT
C2835757|T037|S24.101D|ICD10CM|UNSPECIFIED INJURY AT T1 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY AT T1 LEVEL OF THORACIC SPINAL CORD, SUBS ENCNTR
C2889292|T047|M05.571|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT ANK/FT
C2884036|T037|T51.3X2A|ICD10CM|TOXIC EFFECT OF FUSEL OIL, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF FUSEL OIL, INTENTIONAL SELF-HARM, INIT
C2890260|T037|T83.120A|ICD10CM|DISPLACEMENT OF URINARY ELECTRONIC STIMULATOR DEVICE, INITIAL ENCOUNTER|DISPLACEMENT OF URINARY ELECTRONIC STIMULATOR DEVICE, INIT
C2874245|T047|E71.39|ICD10CM|OTHER DISORDERS OF FATTY-ACID METABOLISM|OTHER DISORDERS OF FATTY-ACID METABOLISM
C2889229|T047|M05.39|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS MULT SITE
C4270607|T046|T85.810A|ICD10CM|EMBOLISM DUE TO NERVOUS SYSTEM PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|EMBOLISM DUE TO NERVOUS SYSTEM PROSTH DEV/GRFT, INIT
C2889198|T047|M05.30|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP SITE
C0268634|T047|E71.30|ICD10CM|DISORDER OF FATTY-ACID METABOLISM, UNSPECIFIED|DISORDER OF FATTY-ACID METABOLISM, UNSPECIFIED
C2874244|T047||ICD10CM|DISORDERS OF KETONE METABOLISM
C2834049|T037|S14.155D|ICD10CM|OTHER INCOMPLETE LESION AT C5 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|OTH INCOMPLETE LESION AT C5, SUBS
C2858612|T037|S72.435C|ICD10CM|NONDISPLACED FRACTURE OF MEDIAL CONDYLE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF MED CONDYLE OF L FEMR, 7THC
C2858611|T037|S72.435B|ICD10CM|NONDISPLACED FRACTURE OF MEDIAL CONDYLE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF MED CONDYLE OF L FEMR, 7THB
C2858610|T037|S72.435A|ICD10CM|NONDISPLACED FRACTURE OF MEDIAL CONDYLE OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF MEDIAL CONDYLE OF LEFT FEMUR, INIT FOR CLOS FX
C2834048|T037|S14.155A|ICD10CM|OTHER INCOMPLETE LESION AT C5 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|OTH INCOMPLETE LESION AT C5, INIT
C2837875|T037|S32.392A|ICD10CM|OTHER FRACTURE OF LEFT ILIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF LEFT ILIUM, INIT ENCNTR FOR CLOSED FRACTURE
C2889330|T047|M05.719|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED SHOULDER WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRIT W RHEU FACTOR OF UNSP SHLDR W/O ORG/SYS INVOLV
C2834050|T037|S14.155S|ICD10CM|OTHER INCOMPLETE LESION AT C5 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|OTH INCOMPLETE LESION AT C5, SEQUELA
C2889329|T047|M05.712|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT SHOULDER WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRIT W RHEU FACTOR OF L SHOULDER W/O ORG/SYS INVOLV
C2889328|T047|M05.711|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT SHOULDER WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRIT W RHEU FACTOR OF R SHOULDER W/O ORG/SYS INVOLV
C2834003|T037|S14.143S|ICD10CM|BROWN-SEQUARD SYNDROME AT C3 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|BROWN-SEQUARD SYNDROME AT C3, SEQUELA
C2865557|T037|S88.121S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, RIGHT LOWER LEG, SEQUELA|PART TRAUM AMP AT LEVEL BETW KNEE AND ANKLE, R LOW LEG, SQLA
C2887762|T047|K50.10|ICD10CM|CROHN'S DISEASE OF LARGE INTESTINE WITHOUT COMPLICATIONS|CROHN'S DISEASE OF LARGE INTESTINE WITHOUT COMPLICATIONS
C2834001|T037|S14.143A|ICD10CM|BROWN-SEQUARD SYNDROME AT C3 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|BROWN-SEQUARD SYNDROME AT C3, INIT
C2834002|T037|S14.143D|ICD10CM|BROWN-SEQUARD SYNDROME AT C3 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|BROWN-SEQUARD SYNDROME AT C3, SUBS
C2884038|T037|T51.3X2S|ICD10CM|TOXIC EFFECT OF FUSEL OIL, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF FUSEL OIL, INTENTIONAL SELF-HARM, SEQUELA
C2875147|T047|G43.011|ICD10CM|MIGRAINE WITHOUT AURA, INTRACTABLE, WITH STATUS MIGRAINOSUS|MIGRAINE WITHOUT AURA, INTRACTABLE, WITH STATUS MIGRAINOSUS
C2875148|T047|G43.019|ICD10CM|MIGRAINE WITHOUT AURA, INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|MIGRAINE W/O AURA, INTRACTABLE, WITHOUT STATUS MIGRAINOSUS
C2833891|T037|S14.113D|ICD10CM|COMPLETE LESION AT C3 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION AT C3 LEVEL OF CERVICAL SPINAL CORD, SUBS
C2884368|T037|T54.1X2S|ICD10CM|TOXIC EFFECT OF OTHER CORROSIVE ORGANIC COMPOUNDS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CORROSIVE ORGANIC COMPND, SELF-HARM, SEQUELA
C2889915|T037|T82.320A|ICD10CM|DISPLACEMENT OF AORTIC (BIFURCATION) GRAFT (REPLACEMENT), INITIAL ENCOUNTER|DISPLACEMENT OF AORTIC (BIFURCATION) GRAFT, INIT
C4268050|T047|E10.3541|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, RIGHT EYE|TYPE 1 DIAB WITH PROLIF DIAB RTNOP WITH COMB DETACH, R EYE
C4268052|T047|E10.3543|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, BILATERAL|TYPE 1 DIAB WITH PROLIF DIABETIC RTNOP WITH COMB DETACH, BI
C4268051|T047|E10.3542|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, LEFT EYE|TYPE 1 DIAB WITH PROLIF DIAB RTNOP WITH COMB DETACH, L EYE
C2887802|T047|K51.218|ICD10CM|ULCERATIVE (CHRONIC) PROCTITIS WITH OTHER COMPLICATION|ULCERATIVE (CHRONIC) PROCTITIS WITH OTHER COMPLICATION
C2887803|T047|K51.219|ICD10CM|ULCERATIVE (CHRONIC) PROCTITIS WITH UNSPECIFIED COMPLICATIONS|ULCERATIVE (CHRONIC) PROCTITIS WITH UNSP COMPLICATIONS
C2887801|T047|K51.214|ICD10CM|ULCERATIVE (CHRONIC) PROCTITIS WITH ABSCESS|ULCERATIVE (CHRONIC) PROCTITIS WITH ABSCESS
C2887798|T047|K51.211|ICD10CM|ULCERATIVE (CHRONIC) PROCTITIS WITH RECTAL BLEEDING|ULCERATIVE (CHRONIC) PROCTITIS WITH RECTAL BLEEDING
C2887799|T047|K51.212|ICD10CM|ULCERATIVE (CHRONIC) PROCTITIS WITH INTESTINAL OBSTRUCTION|ULCERATIVE (CHRONIC) PROCTITIS WITH INTESTINAL OBSTRUCTION
C2887800|T047|K51.213|ICD10CM|ULCERATIVE (CHRONIC) PROCTITIS WITH FISTULA|ULCERATIVE (CHRONIC) PROCTITIS WITH FISTULA
C2833405|T037|S12.331A|ICD10CM|UNSPECIFIED TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP TRAUM NONDISP SPONDYLOLYSIS OF 4TH CERVCAL VERT, INIT
C2833406|T037|S12.331B|ICD10CM|UNSPECIFIED TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP TRAUM NONDISP SPONDYLOLYSIS OF 4TH CERVCAL VERT, 7THB
C2890670|T037|T84.193A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTERNAL FIXATION DEVICE OF BONE OF LEFT FOREARM, INITIAL ENCOUNTER|MECH COMPL OF INT FIX OF BONE OF LEFT FOREARM, INIT
C2838343|T037|S32.486A|ICD10CM|NONDISPLACED DOME FRACTURE OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED DOME FRACTURE OF UNSP ACETABULUM, INIT
C2901032|T046|M84.462A|ICD10CM|PATHOLOGICAL FRACTURE, LEFT TIBIA, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, LEFT TIBIA, INIT ENCNTR FOR FRACTURE
C2837509|T037|S32.019A|ICD10CM|UNSPECIFIED FRACTURE OF FIRST LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF FIRST LUMBAR VERTEBRA, INIT FOR CLOS FX
C2837510|T037|S32.019B|ICD10CM|UNSPECIFIED FRACTURE OF FIRST LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF FIRST LUMBAR VERTEBRA, INIT FOR OPN FX
C2901546|T046|M84.671A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, RIGHT ANKLE, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, RIGHT ANKLE, INIT
C2878686|T037|T43.8X2A|ICD10CM|POISONING BY OTHER PSYCHOTROPIC DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH PSYCHOTROPIC DRUGS, SELF-HARM, INIT
C2887461|T047|J45.51|ICD10CM|SEVERE PERSISTENT ASTHMA WITH (ACUTE) EXACERBATION|SEVERE PERSISTENT ASTHMA WITH (ACUTE) EXACERBATION
C2887460|T047||ICD10CM|SEVERE PERSISTENT ASTHMA, UNCOMPLICATED
C2887462|T047||ICD10CM|SEVERE PERSISTENT ASTHMA WITH STATUS ASTHMATICUS
C2901263|T046|M84.553A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, UNSP FEMUR, INIT
C2838443|T037|S32.613A|ICD10CM|DISPLACED AVULSION FRACTURE OF UNSPECIFIED ISCHIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED AVULSION FRACTURE OF UNSP ISCHIUM, INIT
C2878688|T037|T43.8X2S|ICD10CM|POISONING BY OTHER PSYCHOTROPIC DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH PSYCHOTROPIC DRUGS, SELF-HARM, SEQUELA
C2838444|T037|S32.613B|ICD10CM|DISPLACED AVULSION FRACTURE OF UNSPECIFIED ISCHIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISPLACED AVULSION FRACTURE OF UNSP ISCHIUM, INIT FOR OPN FX
C2874703|T048|F16.288|ICD10CM|HALLUCINOGEN DEPENDENCE WITH OTHER HALLUCINOGEN-INDUCED DISORDER|HALLUCINOGEN DEPENDENCE W OTH HALLUCINOGEN-INDUCED DISORDER
C0582499|T191|C48.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF RETROPERITONEUM AND PERITONEUM|BOESARTIGE NEUBILDUNG: RETROPERITONEUM UND PERITONEUM, MEHRERE TEILBEREICHE UEBERLAPPEND
C2833773|T037|S14.0XXS|ICD10CM|CONCUSSION AND EDEMA OF CERVICAL SPINAL CORD, SEQUELA|CONCUSSION AND EDEMA OF CERVICAL SPINAL CORD, SEQUELA
C2874704|T048|F16.280|ICD10CM|HALLUCINOGEN DEPENDENCE WITH HALLUCINOGEN-INDUCED ANXIETY DISORDER|HALLUCINOGEN DEPENDENCE W ANXIETY DISORDER
C2874705|T048|F16.283|ICD10CM|HALLUCINOGEN DEPENDENCE WITH HALLUCINOGEN PERSISTING PERCEPTION DISORDER (FLASHBACKS)|HALLUCIGN DEPEND W HALLUCIGN PERSISTING PERCEPTION DISORDER
C2890534|T037|T84.061A|ICD10CM|WEAR OF ARTICULAR BEARING SURFACE OF INTERNAL PROSTHETIC LEFT HIP JOINT, INITIAL ENCOUNTER|WEAR OF ARTIC BEARING SURFACE OF INT PROSTH L HIP JT, INIT
C2888922|T047|M00.871|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, RIGHT ANKLE AND FOOT|ARTHRITIS DUE TO OTHER BACTERIA, RIGHT ANKLE AND FOOT
C2888923|T047|M00.872|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, LEFT ANKLE AND FOOT|ARTHRITIS DUE TO OTHER BACTERIA, LEFT ANKLE AND FOOT
C2888924|T047|M00.879|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, UNSPECIFIED ANKLE AND FOOT|ARTHRITIS DUE TO OTHER BACTERIA, UNSPECIFIED ANKLE AND FOOT
C2833771|T037|S14.0XXA|ICD10CM|CONCUSSION AND EDEMA OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|CONCUSSION AND EDEMA OF CERVICAL SPINAL CORD, INIT ENCNTR
C2845939|T191|C72.59|ICD10CM|MALIGNANT NEOPLASM OF OTHER CRANIAL NERVES|MALIGNANT NEOPLASM OF OTHER CRANIAL NERVES
C2833772|T037|S14.0XXD|ICD10CM|CONCUSSION AND EDEMA OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|CONCUSSION AND EDEMA OF CERVICAL SPINAL CORD, SUBS ENCNTR
C4509273|T047|L89.019|ICD10CM|PRESSURE ULCER OF RIGHT ELBOW, UNSPECIFIED STAGE|HEALING PRESSURE ULCER OF RIGHT ELBOW, UNSPECIFIED STAGE
C2888226|T047|L89.012|ICD10CM|PRESSURE ULCER OF RIGHT ELBOW, STAGE 2|PRESSURE ULCER OF RIGHT ELBOW, STAGE 2
C2888229|T047|L89.013|ICD10CM|PRESSURE ULCER OF RIGHT ELBOW, STAGE 3|PRESSURE ULCER OF RIGHT ELBOW, STAGE 3
C2888220|T047||ICD10CM|PRESSURE ULCER OF RIGHT ELBOW, UNSTAGEABLE
C2888223|T047|L89.011|ICD10CM|PRESSURE ULCER OF RIGHT ELBOW, STAGE 1|PRESSURE ULCER OF RIGHT ELBOW, STAGE 1
C2888232|T047|L89.014|ICD10CM|PRESSURE ULCER OF RIGHT ELBOW, STAGE 4|PRESSURE ULCER OF RIGHT ELBOW, STAGE 4
C2882936|T047|I70.631|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF THIGH|ATHSCL NONBIOL BYPASS OF THE RIGHT LEG W ULCERATION OF THIGH
C2882938|T047|I70.633|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF ANKLE|ATHSCL NONBIOL BYPASS OF THE RIGHT LEG W ULCERATION OF ANKLE
C2882937|T047|I70.632|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF CALF|ATHSCL NONBIOL BYPASS OF THE RIGHT LEG W ULCERATION OF CALF
C2882942|T047|I70.635|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF OTHER PART OF FOOT|ATHSCL NONBIOL BYPASS OF THE RIGHT LEG W ULCER OTH PRT FOOT
C2882940|T047|I70.634|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF HEEL AND MIDFOOT|ATHSCL NONBIOL BYPASS OF RIGHT LEG W ULCER OF HEEL AND MIDFT
C2882944|T047|I70.639|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF UNSPECIFIED SITE|ATHSCL NONBIOL BYPASS OF THE RIGHT LEG W ULCER OF UNSP SITE
C2882943|T047|I70.638|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE RIGHT LEG WITH ULCERATION OF OTHER PART OF LOWER LEG|ATHSCL NONBIOL BYPASS OF RIGHT LEG W ULCER OTH PRT LOW LEG
C2838071|T037|S32.424A|ICD10CM|NONDISPLACED FRACTURE OF POSTERIOR WALL OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF POSTERIOR WALL OF RIGHT ACETABULUM, INIT
C2896676|T046|M80.819A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, UNSPECIFIED SHOULDER, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, UNSP SHOULDER, INIT
C2901124|T046|M84.48XA|ICD10CM|PATHOLOGICAL FRACTURE, OTHER SITE, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, OTHER SITE, INIT ENCNTR FOR FRACTURE
C2905727|T037|X77.0XXD|ICD10CM|INTENTIONAL SELF-HARM BY STEAM OR HOT VAPORS, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY STEAM OR HOT VAPORS, SUBS ENCNTR
C2838380|T037|S32.511B|ICD10CM|FRACTURE OF SUPERIOR RIM OF RIGHT PUBIS, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF SUPERIOR RIM OF RIGHT PUBIS, INIT FOR OPN FX
C4509330|T047|L97.906|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF UNSPECIFIED LOWER LEG WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC UNSP PRT UNSP LW LEG W BNE INVL W/O EVD NECR
C4509329|T047|L97.905|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF UNSPECIFIED LOWER LEG WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC UNSP PRT UNSP LW LEG W MSL INVL W/O EVD NECR
C2888758|T047|L97.904|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF UNSPECIFIED LOWER LEG WITH NECROSIS OF BONE|NON-PRS CHRONIC ULC UNSP PRT OF UNSP LOWER LEG W NECROS BONE
C2888757|T047|L97.903|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF UNSPECIFIED LOWER LEG WITH NECROSIS OF MUSCLE|NON-PRS CHRONIC ULC UNSP PRT OF UNSP LOW LEG W NECROS MUSCLE
C2888756|T047|L97.902|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF UNSPECIFIED LOWER LEG WITH FAT LAYER EXPOSED|NON-PRS CHR ULC UNSP PRT OF UNSP LOW LEG W FAT LAYER EXPOSED
C2888755|T047|L97.901|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF UNSPECIFIED LOWER LEG LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHR ULC UNSP PRT OF UNSP LOW LEG LMT TO BRKDWN SKIN
C2901889|T047|M86.479|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, UNSPECIFIED ANKLE AND FOOT|CHRONIC OSTEOMYELITIS W DRAINING SINUS, UNSP ANKLE AND FOOT
C2901888|T047|M86.472|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, LEFT ANKLE AND FOOT|CHRONIC OSTEOMYELITIS W DRAINING SINUS, LEFT ANKLE AND FOOT
C2888759|T047|L97.909|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF UNSPECIFIED LOWER LEG WITH UNSPECIFIED SEVERITY|NON-PRS CHRONIC ULC UNSP PRT OF UNSP LOW LEG W UNSP SEVERITY
C4509331|T047|L97.908|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED PART OF UNSPECIFIED LOWER LEG WITH OTHER SPECIFIED SEVERITY|NON-PRS CHRONIC ULC UNSP PRT OF UNSP LOW LEG WITH OTH SEVERT
C2901212|T046|M84.539A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, UNSPECIFIED ULNA AND RADIUS, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLTC DISEASE, UNSP ULNA AND RADIUS, INIT
C2832678|T037|S06.9X1S|ICD10CM|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|UNSP INTCRN INJURY W LOC OF 30 MINUTES OR LESS, SEQUELA
C2910020|T047|P36.39|ICD10CM|SEPSIS OF NEWBORN DUE TO OTHER STAPHYLOCOCCI|SEPSIS OF NEWBORN DUE TO OTHER STAPHYLOCOCCI
C2858816|T037|S72.455A|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP SUPRCNDL FX W/O INTRCNDL EXTN LOWER END L FEMR, INIT
C2910019|T047|P36.30|ICD10CM|SEPSIS OF NEWBORN DUE TO UNSPECIFIED STAPHYLOCOCCI|SEPSIS OF NEWBORN DUE TO UNSPECIFIED STAPHYLOCOCCI
C2833145|T037|S12.001A|ICD10CM|UNSPECIFIED NONDISPLACED FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP NONDISP FX OF FIRST CERVICAL VERTEBRA, INIT FOR CLOS FX
C2858818|T037|S72.455C|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP SUPRCNDL FX W/O INTRCNDL EXTN LOW END L FEMR, 7THC
C4509245|T047|I50.84|ICD10CM|END STAGE HEART FAILURE|STAGE D HEART FAILURE
C0221045|T047|I50.83|ICD10CM|HIGH OUTPUT HEART FAILURE|HIGH OUTPUT HEART FAILURE
C0685095|T047|I50.82|ICD10CM|BIVENTRICULAR HEART FAILURE|BIVENTRICULAR HEART FAILURE
C2874781|T048|F18.951|ICD10CM|INHALANT USE, UNSPECIFIED WITH INHALANT-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|INHALANT USE, UNSP W INHALNT-INDUCE PSYCH DISORD W HALLUCIN
C2874780|T048|F18.950|ICD10CM|INHALANT USE, UNSPECIFIED WITH INHALANT-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|INHALANT USE, UNSP W INHALNT-INDUCE PSYCH DISORD W DELUSIONS
C2890938|T037|T85.03XA|ICD10CM|LEAKAGE OF VENTRICULAR INTRACRANIAL (COMMUNICATING) SHUNT, INITIAL ENCOUNTER|LEAKAGE OF VENTRICULAR INTRACRANIAL SHUNT, INIT
C2874782|T048|F18.959|ICD10CM|INHALANT USE, UNSPECIFIED WITH INHALANT-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|INHALANT USE, UNSP W INHALNT-INDUCE PSYCHOTIC DISORDER, UNSP
C2901915|T047|M86.61|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, UNSPECIFIED SHOULDER|OTHER CHRONIC OSTEOMYELITIS, SHOULDER
C4268479|T046|I63.213|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF BILATERAL VERTEBRAL ARTERIES|CEREB INFRC DUE TO UNSP OCCLS OR STENOSIS OF BI VERTEB ART
C2882354|T046|I63.212|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF LEFT VERTEBRAL ARTERY|CEREBRAL INFRC DUE TO UNSP OCCLS OR STENOSIS OF L VERTEB ART
C2882353|T046|I63.211|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF RIGHT VERTEBRAL ARTERY|CEREBRAL INFRC DUE TO UNSP OCCLS OR STENOSIS OF R VERTEB ART
C0392096|T033|Z94.0|DMDICD10|KIDNEY TRANSPLANT STATUS|ZUSTAND NACH NIERENTRANSPLANTATION
C2901914|T047|M86.612|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, LEFT SHOULDER|OTHER CHRONIC OSTEOMYELITIS, LEFT SHOULDER
C2838621|T037|S34.102D|ICD10CM|UNSPECIFIED INJURY TO L2 LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY TO L2 LEVEL OF LUMBAR SPINAL CORD, SUBS ENCNTR
C2901913|T047|M86.611|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, RIGHT SHOULDER|OTHER CHRONIC OSTEOMYELITIS, RIGHT SHOULDER
C2882355|T046|I63.219|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF UNSPECIFIED VERTEBRAL ARTERIES|CEREB INFRC DUE TO UNSP OCCLS OR STENOSIS OF UNSP VERTEB ART
C2873995|T047|E09.59|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH OTHER CIRCULATORY COMPLICATIONS|DRUG/CHEM DIABETES MELLITUS W OTH CIRCULATORY COMPLICATIONS
C2842150|T191|C57.02|ICD10CM|MALIGNANT NEOPLASM OF LEFT FALLOPIAN TUBE|MALIGNANT NEOPLASM OF LEFT FALLOPIAN TUBE
C2842148|T191|C57.00|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED FALLOPIAN TUBE|MALIGNANT NEOPLASM OF UNSPECIFIED FALLOPIAN TUBE
C2842149|T191|C57.01|ICD10CM|MALIGNANT NEOPLASM OF RIGHT FALLOPIAN TUBE|MALIGNANT NEOPLASM OF RIGHT FALLOPIAN TUBE
C2905732|T037|X77.1XXS|ICD10CM|INTENTIONAL SELF-HARM BY HOT TAP WATER, SEQUELA|INTENTIONAL SELF-HARM BY HOT TAP WATER, SEQUELA
C3264498|T047|M86.669|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, UNSPECIFIED TIBIA AND FIBULA|OTHER CHRONIC OSTEOMYELITIS, UNSPECIFIED TIBIA AND FIBULA
C2905730|T037|X77.1XXA|ICD10CM|INTENTIONAL SELF-HARM BY HOT TAP WATER, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY HOT TAP WATER, INITIAL ENCOUNTER
C2905731|T037|X77.1XXD|ICD10CM|INTENTIONAL SELF-HARM BY HOT TAP WATER, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY HOT TAP WATER, SUBSEQUENT ENCOUNTER
C2890271|T037|T83.128A|ICD10CM|DISPLACEMENT OF OTHER URINARY DEVICES AND IMPLANTS, INITIAL ENCOUNTER|DISPLACEMENT OF OTH URINARY DEVICES AND IMPLANTS, INIT
C2860089|T037|S79.019A|ICD10CM|SALTER-HARRIS TYPE I PHYSEAL FRACTURE OF UPPER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SLTR-HARIS TYPE I PHYSEAL FX UPPER END OF UNSP FEMUR, INIT
C2832495|T037|S06.5X6S|ICD10CM|TRAUMATIC SUBDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|TRAUM SUBDR HEM W LOC >24 HR W/O RET CONSC W SURV, SEQUELA
C2884152|T037|T52.4X2A|ICD10CM|TOXIC EFFECT OF KETONES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF KETONES, INTENTIONAL SELF-HARM, INIT ENCNTR
C4268298|T048|F19.288|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH OTHER PSYCHOACTIVE SUBSTANCE-INDUCED DISORDER|OTHER (OR UNKNOWN) SUBSTANCE USE DISORDER, SEVERE, WITH OTHER (OR UNKNOWN) SUBSTANCE INDUCED OBSESSIVE-COMPULSIVE OR RELATED DISORDER
C2874828|T048|F19.280|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH PSYCHOACTIVE SUBSTANCE-INDUCED ANXIETY DISORDER|OTH PSYCHOACTIVE SUBSTANCE DEPENDENCE W ANXIETY DISORDER
C2874829|T048|F19.281|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH PSYCHOACTIVE SUBSTANCE-INDUCED SEXUAL DYSFUNCTION|OTH PSYCHOACTIVE SUBSTANCE DEPENDENCE W SEXUAL DYSFUNCTION
C2874830|T048|F19.282|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH PSYCHOACTIVE SUBSTANCE-INDUCED SLEEP DISORDER|OTH PSYCHOACTIVE SUBSTANCE DEPENDENCE W SLEEP DISORDER
C2832493|T037|S06.5X6A|ICD10CM|TRAUMATIC SUBDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|TRAUM SUBDR HEM W LOC >24 HR W/O RET CONSC W SURV, INIT
C2884154|T037|T52.4X2S|ICD10CM|TOXIC EFFECT OF KETONES, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF KETONES, INTENTIONAL SELF-HARM, SEQUELA
C2521520|T060|C01|ICD10PCS|MALIGNANT NEOPLASM OF BASE OF TONGUE|NUCLEAR MEDICINE, CENTRAL NERVOUS SYS, PLANAR NUCL MED IMAG
C0747273|T191|C07|DMDICD10|MALIGNANT NEOPLASM OF PAROTID GLAND|BOESARTIGE NEUBILDUNG DER PAROTIS
C2838622|T037|S34.102S|ICD10CM|UNSPECIFIED INJURY TO L2 LEVEL OF LUMBAR SPINAL CORD, SEQUELA|UNSP INJURY TO L2 LEVEL OF LUMBAR SPINAL CORD, SEQUELA
C2832232|T037|S06.343A|ICD10CM|TRAUMATIC HEMORRHAGE OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 1 HOURS TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|TRAUM HEMOR RIGHT CEREBRUM W LOC OF 1-5 HRS 59 MINUTES, INIT
C2865520|T037|S88.012A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT KNEE LEVEL, LEFT LOWER LEG, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION AT KNEE LEVEL, L LOW LEG, INIT
C2835766|T037|S24.103S|ICD10CM|UNSPECIFIED INJURY AT T7-T10 LEVEL OF THORACIC SPINAL CORD, SEQUELA|UNSP INJURY AT T7-T10 LEVEL OF THORACIC SPINAL CORD, SEQUELA
C2911490|T033|Z93.52|ICD10CM|APPENDICO-VESICOSTOMY STATUS|APPENDICO-VESICOSTOMY STATUS
C2865521|T037|S88.012D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT KNEE LEVEL, LEFT LOWER LEG, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION AT KNEE LEVEL, L LOW LEG, SUBS
C2832234|T037|S06.343S|ICD10CM|TRAUMATIC HEMORRHAGE OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 1 HOURS TO 5 HOURS 59 MINUTES, SEQUELA|TRAUM HEMOR R CEREB W LOC OF 1-5 HRS 59 MINUTES, SEQUELA
C2865522|T037|S88.012S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT KNEE LEVEL, LEFT LOWER LEG, SEQUELA|COMPLETE TRAUMATIC AMP AT KNEE LEVEL, L LOW LEG, SEQUELA
C2833637|T037|S12.690B|ICD10CM|OTHER DISPLACED FRACTURE OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH DISP FX OF SEVENTH CERVICAL VERTEBRA, INIT FOR OPN FX
C2838686|T037|S34.129A|ICD10CM|INCOMPLETE LESION OF UNSPECIFIED LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|INCOMPLETE LESION OF UNSP LEVEL OF LUMBAR SPINAL CORD, INIT
C2833636|T037|S12.690A|ICD10CM|OTHER DISPLACED FRACTURE OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH DISP FX OF SEVENTH CERVICAL VERTEBRA, INIT FOR CLOS FX
C4268091|T047|E11.3499|ICD10CM|TYPE 2 DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|TYPE 2 DIAB WITH SEVERE NONP RTNOP WITHOUT MCLR EDEMA, UNSP
C4268089|T047|E11.3492|ICD10CM|TYPE 2 DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|TYPE 2 DIAB WITH SEVERE NONP RTNOP WITHOUT MCLR EDEMA, L EYE
C4268090|T047|E11.3493|ICD10CM|TYPE 2 DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|TYPE 2 DIAB WITH SEVERE NONP RTNOP WITHOUT MACULAR EDEMA, BI
C4268088|T047|E11.3491|ICD10CM|TYPE 2 DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|TYPE 2 DIAB WITH SEVERE NONP RTNOP WITHOUT MCLR EDEMA, R EYE
C2856568|T037|S72.019A|ICD10CM|UNSPECIFIED INTRACAPSULAR FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP INTRACAPSULAR FRACTURE OF UNSP FEMUR, INIT FOR CLOS FX
C2856570|T037|S72.019C|ICD10CM|UNSPECIFIED INTRACAPSULAR FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP INTRACAP FX UNSP FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2875177|T047|G43.719|ICD10CM|CHRONIC MIGRAINE WITHOUT AURA, INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|CHRONIC MIGRAINE W/O AURA, INTRACTABLE, W/O STAT MIGR
C2875176|T047|G43.711|ICD10CM|CHRONIC MIGRAINE WITHOUT AURA, INTRACTABLE, WITH STATUS MIGRAINOSUS|CHRONIC MIGRAINE W/O AURA, INTRACTABLE, W STATUS MIGRAINOSUS
C2890902|T037|T84.82XA|ICD10CM|FIBROSIS DUE TO INTERNAL ORTHOPEDIC PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|FIBROSIS DUE TO INTERNAL ORTHOPEDIC PROSTH DEV/GRFT, INIT
C2832575|T037|S06.816S|ICD10CM|INJURY OF RIGHT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|INJ R INT CRTD,INTCR W LOC >24 HR W/O RET CONSC W SURV, SQLA
C2888889|T047|M00.272|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, LEFT ANKLE AND FOOT|OTHER STREPTOCOCCAL ARTHRITIS, LEFT ANKLE AND FOOT
C2874760|T048||ICD10CM|INHALANT DEPENDENCE WITH INTOXICATION, UNCOMPLICATED
C2888888|T047|M00.271|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, RIGHT ANKLE AND FOOT|OTHER STREPTOCOCCAL ARTHRITIS, RIGHT ANKLE AND FOOT
C2873984|T047|E09.41|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH NEUROLOGICAL COMPLICATIONS WITH DIABETIC MONONEUROPATHY|DRUG/CHEM DIABETES W NEURO COMP W DIABETIC MONONEUROPATHY
C2874762|T048|F18.229|ICD10CM|INHALANT DEPENDENCE WITH INTOXICATION, UNSPECIFIED|INHALANT DEPENDENCE WITH INTOXICATION, UNSPECIFIED
C2835786|T037|S24.113S|ICD10CM|COMPLETE LESION AT T7-T10 LEVEL OF THORACIC SPINAL CORD, SEQUELA|COMPLETE LESION AT T7-T10, SEQUELA
C2888890|T047|M00.279|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, UNSPECIFIED ANKLE AND FOOT|OTHER STREPTOCOCCAL ARTHRITIS, UNSPECIFIED ANKLE AND FOOT
C2832573|T037|S06.816A|ICD10CM|INJURY OF RIGHT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|INJ R INT CRTD,INTCR W LOC >24 HR W/O RET CONSC W SURV, INIT
C2873988|T047|E09.43|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH NEUROLOGICAL COMPLICATIONS WITH DIABETIC AUTONOMIC (POLY)NEUROPATHY|DRUG/CHEM DIAB W NEURO COMP W DIAB AUTONM (POLY)NEUROPATHY
C0837437|T047|M02.30|ICD10AM|REITER'S DISEASE, UNSPECIFIED SITE|REITER'S DISEASE, MULTIPLE SITES
C2873986|T047|E09.42|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH NEUROLOGICAL COMPLICATIONS WITH DIABETIC POLYNEUROPATHY|DRUG/CHEM DIABETES W NEUROLOGICAL COMP W DIABETIC POLYNEUROP
C0837437|T047|M02.39|ICD10CM|REITER'S DISEASE, MULTIPLE SITES|REITER'S DISEASE, MULTIPLE SITES
C2889077|T047|M02.38|ICD10CM|REITER'S DISEASE, VERTEBRAE|REITER'S DISEASE, VERTEBRAE
C2832455|T037|S06.4X6S|ICD10CM|EPIDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|EPIDURAL HEMOR W LOC >24 HR W/O RET CONSC W SURV, SEQUELA
C2889546|T047|M08.071|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, RIGHT ANKLE AND FOOT|UNSP JUVENILE RHEUMATOID ARTHRITIS, RIGHT ANKLE AND FOOT
C2889547|T047|M08.072|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, LEFT ANKLE AND FOOT|UNSP JUVENILE RHEUMATOID ARTHRITIS, LEFT ANKLE AND FOOT
C2889548|T047|M08.079|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED ANKLE AND FOOT|UNSP JUVENILE RHEUMATOID ARTHRITIS, UNSP ANKLE AND FOOT
C2890087|T037|T82.538A|ICD10CM|LEAKAGE OF OTHER CARDIAC AND VASCULAR DEVICES AND IMPLANTS, INITIAL ENCOUNTER|LEAKAGE OF CARDIAC AND VASCULAR DEVICES AND IMPLANTS, INIT
C2905795|T037|X82.1XXD|ICD10CM|INTENTIONAL COLLISION OF MOTOR VEHICLE WITH TRAIN, SUBSEQUENT ENCOUNTER|INTENTIONAL COLLISION OF MOTOR VEHICLE W TRAIN, SUBS ENCNTR
C4270270|T046|T83.192A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INDWELLING URETERAL STENT, INITIAL ENCOUNTER|MECH COMPL OF INDWELLING URETERAL STENT, INITIAL ENCOUNTER
C2857121|T037|S72.102B|ICD10CM|UNSPECIFIED TROCHANTERIC FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP TROCHAN FX LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C2857122|T037|S72.102C|ICD10CM|UNSPECIFIED TROCHANTERIC FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP TROCHAN FX LEFT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2857120|T037|S72.102A|ICD10CM|UNSPECIFIED TROCHANTERIC FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP TROCHANTERIC FRACTURE OF LEFT FEMUR, INIT FOR CLOS FX
C4270144|T046|T82.838A|ICD10CM|HEMORRHAGE DUE TO VASCULAR PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|HEMORRHAGE DUE TO VASCULAR PROSTH DEV/GRFT, INIT
C2878202|T037|T42.6X2S|ICD10CM|POISONING BY OTHER ANTIEPILEPTIC AND SEDATIVE-HYPNOTIC DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY OTH ANTIEPLPTC AND SED-HYPNTC DRUGS, SLF-HRM, SQLA
C2888957|T047|M01.X72|ICD10CM|DIRECT INFECTION OF LEFT ANKLE AND FOOT IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIR INFCT OF LEFT ANK/FT IN INFEC/PARASTC DIS CLASSD ELSWHR
C2889118|T047|M05.039|ICD10CM|FELTY'S SYNDROME, UNSPECIFIED WRIST|FELTY'S SYNDROME, UNSPECIFIED WRIST
C2845908|T191|C69.30|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED CHOROID|MALIGNANT NEOPLASM OF UNSPECIFIED CHOROID
C2845909|T191|C69.31|ICD10CM|MALIGNANT NEOPLASM OF RIGHT CHOROID|MALIGNANT NEOPLASM OF RIGHT CHOROID
C2845910|T191|C69.32|ICD10CM|MALIGNANT NEOPLASM OF LEFT CHOROID|MALIGNANT NEOPLASM OF LEFT CHOROID
C2889117|T047|M05.032|ICD10CM|FELTY'S SYNDROME, LEFT WRIST|FELTY'S SYNDROME, LEFT WRIST
C2889116|T047|M05.031|ICD10CM|FELTY'S SYNDROME, RIGHT WRIST|FELTY'S SYNDROME, RIGHT WRIST
C2878200|T037|T42.6X2A|ICD10CM|POISONING BY OTHER ANTIEPILEPTIC AND SEDATIVE-HYPNOTIC DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY OTH ANTIEPLPTC AND SED-HYPNTC DRUGS, SLF-HRM, INIT
C2843316|T037|S48.129A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN UNSPECIFIED SHOULDER AND ELBOW, INITIAL ENCOUNTER|PARTIAL TRAUM AMP AT LEVEL BETW UNSP SHLDR AND ELBOW, INIT
C2889139|T047|M05.121|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT ELBOW|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF R ELBOW
C2879595|T037|T46.8X2S|ICD10CM|POISONING BY ANTIVARICOSE DRUGS, INCLUDING SCLEROSING AGENTS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY ANTIVARIC DRUGS, INC SCLER AGENTS, SLF-HRM, SEQUELA
C4270319|T046|T83.512A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO NEPHROSTOMY CATHETER, INITIAL ENCOUNTER|I/I REACT D/T NEPHROSTOMY CATHETER, INITIAL ENCOUNTER
C2874431|T048|F11.159|ICD10CM|OPIOID ABUSE WITH OPIOID-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|OPIOID ABUSE WITH OPIOID-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED
C2889479|T047|M06.842|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, LEFT HAND|OTHER SPECIFIED RHEUMATOID ARTHRITIS, LEFT HAND
C2837669|T037|S32.110A|ICD10CM|NONDISPLACED ZONE I FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED ZONE I FRACTURE OF SACRUM, INIT FOR CLOS FX
C2837670|T037|S32.110B|ICD10CM|NONDISPLACED ZONE I FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISPLACED ZONE I FRACTURE OF SACRUM, INIT FOR OPN FX
C2874429|T048|F11.150|ICD10CM|OPIOID ABUSE WITH OPIOID-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|OPIOID ABUSE W OPIOID-INDUCED PSYCHOTIC DISORDER W DELUSIONS
C2874430|T048|F11.151|ICD10CM|OPIOID ABUSE WITH OPIOID-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|OPIOID ABUSE W OPIOID-INDUCED PSYCHOTIC DISORDER W HALLUCIN
C2859171|T037|S73.013A|ICD10CM|POSTERIOR SUBLUXATION OF UNSPECIFIED HIP, INITIAL ENCOUNTER|POSTERIOR SUBLUXATION OF UNSPECIFIED HIP, INITIAL ENCOUNTER
C2832150|T037|S06.323S|ICD10CM|CONTUSION AND LACERATION OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, SEQUELA|CONTUS/LAC LEFT CEREBRUM W LOC OF 1-5 HRS 59 MIN, SEQUELA
C0432422|T049|Q91.1|DMDICD10|TRISOMY 18, MOSAICISM (MITOTIC NONDISJUNCTION)|TRISOMIE 18, MOSAIK (MITOTISCHE NON-DISJUNCTION)
C2910354|T047||ICD10CM|TRISOMY 18, NONMOSAICISM (MEIOTIC NONDISJUNCTION)
C3537048|T049|Q91.3|ICD10CM|TRISOMY 18, UNSPECIFIED|TRISOMY 18, UNSPECIFIED
C0432487|T191||ICD10CM|POST-TRANSPLANT LYMPHOPROLIFERATIVE DISORDER (PTLD)
C0017531|T047||ICD10CM|CASTLEMAN DISEASE
C2858113|T037|S72.356A|ICD10CM|NONDISPLACED COMMINUTED FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP COMMINUTED FRACTURE OF SHAFT OF UNSP FEMUR, INIT
C2873721|T191|D47.Z9|ICD10CM|OTHER SPECIFIED NEOPLASMS OF UNCERTAIN BEHAVIOR OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE|HISTIOCYTIC TUMORS OF UNCERTAIN BEHAVIOR
C2858115|T037|S72.356C|ICD10CM|NONDISPLACED COMMINUTED FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP COMMNT FX SHAFT OF UNSP FEMR, 7THC
C2858114|T037|S72.356B|ICD10CM|NONDISPLACED COMMINUTED FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP COMMNT FX SHAFT OF UNSP FEMR, 7THB
C2889692|T037|T81.592D|ICD10CM|OTHER COMPLICATIONS OF FOREIGN BODY ACCIDENTALLY LEFT IN BODY FOLLOWING KIDNEY DIALYSIS, SUBSEQUENT ENCOUNTER|OTH COMP OF FB ACC LEFT IN BODY FOL KIDNEY DIALYSIS, SUBS
C1660761|T047||ICD10CM|PARAPLEGIA, INCOMPLETE
C0030486|T047|G82.2|ICD10CM|PARAPLEGIA, UNSPECIFIED|PARAPLEGIA
C1659098|T047||ICD10CM|PARAPLEGIA, COMPLETE
C2887122|T047|I82.722|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF DEEP VEINS OF LEFT UPPER EXTREMITY|CHRONIC EMBOLISM AND THROMBOSIS OF DEEP VEINS OF L UP EXTREM
C2887123|T047|I82.723|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF DEEP VEINS OF UPPER EXTREMITY, BILATERAL|CHRONIC EMBOLISM AND THOMBOS OF DEEP VEINS OF UP EXTREM, BI
C2887121|T047|I82.721|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF DEEP VEINS OF RIGHT UPPER EXTREMITY|CHRONIC EMBOLISM AND THROMBOSIS OF DEEP VEINS OF R UP EXTREM
C2889693|T037|T81.592S|ICD10CM|OTHER COMPLICATIONS OF FOREIGN BODY ACCIDENTALLY LEFT IN BODY FOLLOWING KIDNEY DIALYSIS, SEQUELA|OTH COMP OF FB ACC LEFT IN BODY FOL KIDNEY DIALYSIS, SEQUELA
C2883560|T037|T50.1X2S|ICD10CM|POISONING BY LOOP [HIGH-CEILING] DIURETICS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY LOOP DIURETICS, INTENTIONAL SELF-HARM, SEQUELA
C2887124|T047|I82.729|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF DEEP VEINS OF UNSPECIFIED UPPER EXTREMITY|CHRONIC EMBOLISM AND THROMBOSIS OF DEEP VN UNSP UP EXTREM
C2902866|T046|N02.0|ICD10CM|RECURRENT AND PERSISTENT HEMATURIA WITH MINOR GLOMERULAR ABNORMALITY|RECURRENT AND PERSISTENT HEMATURIA WITH MINIMAL CHANGE LESION
C2902869|T046|N02.1|ICD10CM|RECURRENT AND PERSISTENT HEMATURIA WITH FOCAL AND SEGMENTAL GLOMERULAR LESIONS|RECURRENT AND PERSISTENT HEMATURIA WITH FOCAL GLOMERULONEPHRITIS
C0475540|T047|N02.2|DMDICD10|RECURRENT AND PERSISTENT HEMATURIA WITH DIFFUSE MEMBRANOUS GLOMERULONEPHRITIS|REZIDIVIERENDE UND PERSISTIERENDE HAEMATURIE: DIFFUSE MEMBRANOESE GLOMERULONEPHRITIS
C0475541|T047|N02.3|DMDICD10|RECURRENT AND PERSISTENT HEMATURIA WITH DIFFUSE MESANGIAL PROLIFERATIVE GLOMERULONEPHRITIS|REZIDIVIERENDE UND PERSISTIERENDE HAEMATURIE: DIFFUSE MESANGIOPROLIFERATIVE GLOMERULONEPHRITIS
C0475542|T047|N02.4|DMDICD10|RECURRENT AND PERSISTENT HEMATURIA WITH DIFFUSE ENDOCAPILLARY PROLIFERATIVE GLOMERULONEPHRITIS|REZIDIVIERENDE UND PERSISTIERENDE HAEMATURIE: DIFFUSE ENDOKAPILLAER-PROLIFERATIVE GLOMERULONEPHRITIS
C2902870|T046|N02.5|ICD10CM|RECURRENT AND PERSISTENT HEMATURIA WITH DIFFUSE MESANGIOCAPILLARY GLOMERULONEPHRITIS|RECURRENT AND PERSISTENT HEMATURIA WITH MEMBRANOPROLIFERATIVE GLOMERULONEPHRITIS, TYPES 1 AND 3, OR NOS
C2896611|T046|M80.069A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, UNSPECIFIED LOWER LEG, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, UNSP LOW LEG, INIT
C2902872|T047|N02.7|ICD10CM|RECURRENT AND PERSISTENT HEMATURIA WITH DIFFUSE CRESCENTIC GLOMERULONEPHRITIS|RECURRENT AND PERSISTENT HEMATURIA WITH EXTRACAPILLARY GLOMERULONEPHRITIS
C2902874|T046|N02.8|ICD10CM|RECURRENT AND PERSISTENT HEMATURIA WITH OTHER MORPHOLOGIC CHANGES|RECURRENT AND PERSISTENT HEMATURIA W OTH MORPHOLOGIC CHANGES
C2902875|T046|N02.9|ICD10CM|RECURRENT AND PERSISTENT HEMATURIA WITH UNSPECIFIED MORPHOLOGIC CHANGES|RECURRENT AND PERST HEMATURIA W UNSP MORPHOLOGIC CHANGES
C2889082|T047|M02.821|ICD10CM|OTHER REACTIVE ARTHROPATHIES, RIGHT ELBOW|OTHER REACTIVE ARTHROPATHIES, RIGHT ELBOW
C2886920|T037|T81.512D|ICD10CM|ADHESIONS DUE TO FOREIGN BODY ACCIDENTALLY LEFT IN BODY FOLLOWING KIDNEY DIALYSIS, SUBSEQUENT ENCOUNTER|ADHES DUE TO FB ACC LEFT IN BODY FOL KIDNEY DIALYSIS, SUBS
C2889083|T047|M02.822|ICD10CM|OTHER REACTIVE ARTHROPATHIES, LEFT ELBOW|OTHER REACTIVE ARTHROPATHIES, LEFT ELBOW
C2886744|T037|T79.8XXA|ICD10CM|OTHER EARLY COMPLICATIONS OF TRAUMA, INITIAL ENCOUNTER|OTHER EARLY COMPLICATIONS OF TRAUMA, INITIAL ENCOUNTER
C2848432|T037|S58.122A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN ELBOW AND WRIST, LEFT ARM, INITIAL ENCOUNTER|PART TRAUM AMP AT LEVEL BETW ELBOW AND WRIST, LEFT ARM, INIT
C2835471|T037|S22.089B|ICD10CM|UNSPECIFIED FRACTURE OF T11-T12 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF T11-T12 VERTEBRA, INIT FOR OPN FX
C2835470|T037|S22.089A|ICD10CM|UNSPECIFIED FRACTURE OF T11-T12 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF T11-T12 VERTEBRA, INIT FOR CLOS FX
C2848434|T037|S58.122S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN ELBOW AND WRIST, LEFT ARM, SEQUELA|PART TRAUM AMP AT LEVEL BETW ELBOW AND WRIST, LEFT ARM, SQLA
C2886364|T037|T71.132A|ICD10CM|ASPHYXIATION DUE TO BEING TRAPPED IN BED LINENS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|ASPHYX DUE TO BEING TRAPPED IN BED LINENS, SELF-HARM, INIT
C4267860|T191|C81.38|ICD10CM|LYMPHOCYTE DEPLETED HODGKIN LYMPHOMA, LYMPH NODES OF MULTIPLE SITES|LYMPHOCYTE DEPLETED HODGKIN LYMPHOMA, LYMPH NODES MULT SITE
C4267861|T191|C81.39|ICD10CM|LYMPHOCYTE DEPLETED HODGKIN LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES|LYMPHOCY DEPLET HODGKIN LYMPH, EXTRNOD AND SOLID ORGAN SITES
C4267854|T191|C81.32|ICD10CM|LYMPHOCYTE DEPLETED HODGKIN LYMPHOMA, INTRATHORACIC LYMPH NODES|LYMPHOCYTE DEPLETED HODGKIN LYMPHOMA, INTRATHORAC NODES
C4267855|T191|C81.33|ICD10CM|LYMPHOCYTE DEPLETED HODGKIN LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES|LYMPHOCYTE DEPLETED HODGKIN LYMPHOMA, INTRA-ABD LYMPH NODES
C4267852|T191|C81.30|ICD10CM|LYMPHOCYTE DEPLETED HODGKIN LYMPHOMA, UNSPECIFIED SITE|LYMPHOCYTE DEPLETED HODGKIN LYMPHOMA, UNSPECIFIED SITE
C4267853|T191|C81.31|ICD10CM|LYMPHOCYTE DEPLETED HODGKIN LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK|LYMPHOCY DEPLET HODGKIN LYMPH, NODES OF HEAD, FACE, AND NECK
C4267858|T191|C81.36|ICD10CM|LYMPHOCYTE DEPLETED HODGKIN LYMPHOMA, INTRAPELVIC LYMPH NODES|LYMPHOCYTE DEPLETED HODGKIN LYMPHOMA, INTRAPELV LYMPH NODES
C4267859|T191|C81.37|ICD10CM|LYMPHOCYTE DEPLETED HODGKIN LYMPHOMA, SPLEEN|LYMPHOCYTE DEPLETED HODGKIN LYMPHOMA, SPLEEN
C4267856|T191|C81.34|ICD10CM|LYMPHOCYTE DEPLETED HODGKIN LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB|LYMPHOCY DEPLET HDGKN LYMPH, NODES OF AXILLA AND UPPER LIMB
C4267857|T191|C81.35|ICD10CM|LYMPHOCYTE DEPLETED HODGKIN LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|LYMPHOCY DEPLET HDGKN LYMPH, NODES OF ING RGN AND LOWER LIMB
C2890794|T037|T84.490A|ICD10CM|OTHER MECHANICAL COMPLICATION OF MUSCLE AND TENDON GRAFT, INITIAL ENCOUNTER|MECH COMPL OF MUSCLE AND TENDON GRAFT, INITIAL ENCOUNTER
C2888999|T047|M02.129|ICD10CM|POSTDYSENTERIC ARTHROPATHY, UNSPECIFIED ELBOW|POSTDYSENTERIC ARTHROPATHY, UNSPECIFIED ELBOW
C2888997|T047|M02.121|ICD10CM|POSTDYSENTERIC ARTHROPATHY, RIGHT ELBOW|POSTDYSENTERIC ARTHROPATHY, RIGHT ELBOW
C2888998|T047|M02.122|ICD10CM|POSTDYSENTERIC ARTHROPATHY, LEFT ELBOW|POSTDYSENTERIC ARTHROPATHY, LEFT ELBOW
C2891271|T037|T86.19|ICD10CM|OTHER COMPLICATION OF KIDNEY TRANSPLANT|OTHER COMPLICATION OF KIDNEY TRANSPLANT
C2891269|T037|T86.10|ICD10CM|UNSPECIFIED COMPLICATION OF KIDNEY TRANSPLANT|UNSPECIFIED COMPLICATION OF KIDNEY TRANSPLANT
C0238217|T046|T86.11|ICD10CM|KIDNEY TRANSPLANT REJECTION|KIDNEY TRANSPLANT REJECTION
C1404117|T046||ICD10CM|KIDNEY TRANSPLANT FAILURE
C2891270|T037|T86.13|ICD10CM|KIDNEY TRANSPLANT INFECTION|KIDNEY TRANSPLANT INFECTION
C4509112|T048|F19.21|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE, IN REMISSION|OTHER (OR UNKNOWN) SUBSTANCE USE, SEVERE, IN SUSTAINED REMISSION
C4237260|T048|F19.20|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE, UNCOMPLICATED|OTHER (OR UNKNOWN) SUBSTANCE USE DISORDER, SEVERE
C0451679|T047|G45.2|DMDICD10|MULTIPLE AND BILATERAL PRECEREBRAL ARTERY SYNDROMES|MULTIPLE UND BILATERALE SYNDROME DER EXTRAZEREBRALEN HIRNVERSORGENDEN ARTERIEN
C2874826|T048|F19.26|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH PSYCHOACTIVE SUBSTANCE-INDUCED PERSISTING AMNESTIC DISORDER|OTH PSYCHOACTV SUBSTANCE DEPEND W PERSIST AMNESTIC DISORDER
C0042568|T047|G45.0|DMDICD10|VERTEBRO-BASILAR ARTERY SYNDROME|ARTERIA-VERTEBRALIS-SYNDROM MIT BASILARIS-SYMPTOMATIK
C0451678|T047|G45.1|DMDICD10|CAROTID ARTERY SYNDROME (HEMISPHERIC)|ARTERIA-CAROTIS-INTERNA-SYNDROM (HALBSEITIG)
C2874832|T048|F19.29|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH UNSPECIFIED PSYCHOACTIVE SUBSTANCE-INDUCED DISORDER|OTH PSYCHOACTIVE SUBSTANCE DEPENDENCE W UNSP DISORDER
C0477375|T047|G45.8|DMDICD10|OTHER TRANSIENT CEREBRAL ISCHEMIC ATTACKS AND RELATED SYNDROMES|SONSTIGE ZEREBRALE TRANSITORISCHE ISCHAEMISCHE ATTACKEN UND VERWANDTE SYNDROME
C0917805|T047||ICD10CM|TRANSIENT CEREBRAL ISCHEMIC ATTACK, UNSPECIFIED
C0348815|T047|E84.0|DMDICD10|CYSTIC FIBROSIS WITH PULMONARY MANIFESTATIONS|ZYSTISCHE FIBROSE MIT LUNGENMANIFESTATIONEN
C0010674|T047|E84.9|DMDICD10|CYSTIC FIBROSIS, UNSPECIFIED|ZYSTISCHE FIBROSE, NICHT NAEHER BEZEICHNET
C0867450|T067|E848|MTHICD9|CYSTIC FIBROSIS WITH OTHER MANIFESTATIONS|ACCIDENT TO, ON, OR INVOLVING, NONMOTOR, NONROAD VEHICLE NOS
C2882200|T047|I25.761|ICD10CM|ATHEROSCLEROSIS OF BYPASS GRAFT OF CORONARY ARTERY OF TRANSPLANTED HEART WITH ANGINA PECTORIS WITH DOCUMENTED SPASM|ATHSCL BYPASS OF COR ART OF TXPLT HEART W ANG PCTRS W SPASM
C2882199|T047|I25.760|ICD10CM|ATHEROSCLEROSIS OF BYPASS GRAFT OF CORONARY ARTERY OF TRANSPLANTED HEART WITH UNSTABLE ANGINA|ATHSCL BYPASS OF COR ART OF TXPLT HEART W UNSTABLE ANGINA
C2882202|T047|I25.769|ICD10CM|ATHEROSCLEROSIS OF BYPASS GRAFT OF CORONARY ARTERY OF TRANSPLANTED HEART WITH UNSPECIFIED ANGINA PECTORIS|ATHSCL BYPASS OF COR ART OF TXPLT HEART W UNSP ANG PCTRS
C2882201|T047|I25.768|ICD10CM|ATHEROSCLEROSIS OF BYPASS GRAFT OF CORONARY ARTERY OF TRANSPLANTED HEART WITH OTHER FORMS OF ANGINA PECTORIS|ATHSCL BYPASS OF COR ART OF TXPLT HEART W OTH ANG PCTRS
C4269280|T037|S02.11AB|ICD10CM|TYPE I OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE I OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, 7THB
C4269279|T037|S02.11AA|ICD10CM|TYPE I OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE I OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, INIT
C4269284|T037|S02.11AS|ICD10CM|TYPE I OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, SEQUELA|TYPE I OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, SEQUELA
C2882591|T047|I69.359|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING CEREBRAL INFARCTION AFFECTING UNSPECIFIED SIDE|HEMIPLGA FOLLOWING CEREBRAL INFARCTION AFFECTING UNSP SIDE
C2882590|T047|I69.354|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING CEREBRAL INFARCTION AFFECTING LEFT NON-DOMINANT SIDE|HEMIPLGA FOLLOWING CEREBRAL INFRC AFFECTING LEFT NONDOM SIDE
C2889966|T037|T82.392A|ICD10CM|OTHER MECHANICAL COMPLICATION OF FEMORAL ARTERIAL GRAFT (BYPASS), INITIAL ENCOUNTER|MECH COMPL OF FEMORAL ARTERIAL GRAFT (BYPASS), INIT ENCNTR
C0869082|T019|Q85.8|DMDICD10|OTHER PHAKOMATOSES, NOT ELSEWHERE CLASSIFIED|SONSTIGE PHAKOMATOSEN, ANDERENORTS NICHT KLASSIFIZIERT
C2882587|T047|I69.351|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING CEREBRAL INFARCTION AFFECTING RIGHT DOMINANT SIDE|HEMIPLGA FOLLOWING CEREBRAL INFRC AFF RIGHT DOMINANT SIDE
C2882588|T047|I69.352|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING CEREBRAL INFARCTION AFFECTING LEFT DOMINANT SIDE|HEMIPLGA FOLLOWING CEREBRAL INFRC AFF LEFT DOMINANT SIDE
C2882589|T047|I69.353|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING CEREBRAL INFARCTION AFFECTING RIGHT NON-DOMINANT SIDE|HEMIPLGA FOLLOWING CEREBRAL INFRC AFF RIGHT NONDOM SIDE
C2896582|T046|M80.052A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, LEFT FEMUR, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, LEFT FEMUR, INIT
C2861603|T191|C92.61|ICD10CM|ACUTE MYELOID LEUKEMIA WITH 11Q23-ABNORMALITY IN REMISSION|ACUTE MYELOID LEUKEMIA WITH 11Q23-ABNORMALITY IN REMISSION
C2861602|T191|C92.60|ICD10CM|ACUTE MYELOID LEUKEMIA WITH 11Q23-ABNORMALITY NOT HAVING ACHIEVED REMISSION|ACUTE MYELOID LEUKEMIA W 11Q23-ABNORMALITY NOT ACHIEVE REMIS
C2861604|T191|C92.62|ICD10CM|ACUTE MYELOID LEUKEMIA WITH 11Q23-ABNORMALITY IN RELAPSE|ACUTE MYELOID LEUKEMIA WITH 11Q23-ABNORMALITY IN RELAPSE
C2838251|T037|S32.465B|ICD10CM|NONDISPLACED ASSOCIATED TRANSVERSE-POSTERIOR FRACTURE OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP ASSOC TRANSV/POST FX LEFT ACETAB, INIT FOR OPN FX
C2838250|T037|S32.465A|ICD10CM|NONDISPLACED ASSOCIATED TRANSVERSE-POSTERIOR FRACTURE OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP ASSOCIATED TRANSV/POST FX LEFT ACETABULUM, INIT
C2888811|T047|M00.049|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, UNSPECIFIED HAND|STAPHYLOCOCCAL ARTHRITIS, UNSPECIFIED HAND
C2833421|T037|S12.350B|ICD10CM|OTHER TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH TRAUM DISPL SPONDYLOLYSIS OF 4TH CERVCAL VERT, 7THB
C2888809|T047|M00.041|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, RIGHT HAND|STAPHYLOCOCCAL ARTHRITIS, RIGHT HAND
C0032463|T191|D45|DMDICD10|POLYCYTHEMIA VERA|POLYCYTHAEMIA VERA
C2888810|T047|M00.042|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, LEFT HAND|STAPHYLOCOCCAL ARTHRITIS, LEFT HAND
C2832032|T037|S06.2X5A|ICD10CM|DIFFUSE TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVELS, INITIAL ENCOUNTER|DIFFUSE TBI W LOC >24 HR W RETURN TO CONSCIOUS LEVELS, INIT
C2832034|T037|S06.2X5S|ICD10CM|DIFFUSE TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVELS, SEQUELA|DIFFUSE TBI W LOC >24 HR W RETURN TO CONSC LEVELS, SEQUELA
C2910104|T019|Q06.9|ICD10CM|CONGENITAL MALFORMATION OF SPINAL CORD, UNSPECIFIED|CONGENITAL DISEASE OR LESION NOS OF SPINAL CORD
C0477975|T019|Q06.8|DMDICD10|OTHER SPECIFIED CONGENITAL MALFORMATIONS OF SPINAL CORD|SONSTIGE NAEHER BEZEICHNETE ANGEBORENE FEHLBILDUNGEN DES RUECKENMARKS
C2833912|T037|S14.118S|ICD10CM|COMPLETE LESION AT C8 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|COMPLETE LESION AT C8 LEVEL OF CERVICAL SPINAL CORD, SEQUELA
C0495480|T019|Q06.1|DMDICD10|HYPOPLASIA AND DYSPLASIA OF SPINAL CORD|HYPOPLASIE UND DYSPLASIE DES RUECKENMARKS
C0266510|T019|Q06.0|DMDICD10|AMYELIA|AMYELIE
C0477974|T019|Q06.3|DMDICD10|OTHER CONGENITAL CAUDA EQUINA MALFORMATIONS|SONSTIGE ANGEBORENE FEHLBILDUNGEN DER CAUDA EQUINA
C0011999|T019|Q06.2|DMDICD10|DIASTEMATOMYELIA|DIASTEMATOMYELIE
C0152444|T047|Q06.4|DMDICD10|HYDROMYELIA|HYDROMYELIE
C2833910|T037|S14.118A|ICD10CM|COMPLETE LESION AT C8 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION AT C8 LEVEL OF CERVICAL SPINAL CORD, INIT
C2833911|T037|S14.118D|ICD10CM|COMPLETE LESION AT C8 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION AT C8 LEVEL OF CERVICAL SPINAL CORD, SUBS
C2859010|T037|S72.499A|ICD10CM|OTHER FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF LOWER END OF UNSP FEMUR, INIT FOR CLOS FX
C2859012|T037|S72.499C|ICD10CM|OTHER FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|OTH FX LOWER END OF UNSP FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2859011|T037|S72.499B|ICD10CM|OTHER FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|OTH FX LOWER END OF UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2877021|T037|T38.1X2A|ICD10CM|POISONING BY THYROID HORMONES AND SUBSTITUTES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY THYROID HORMONES AND SUB, SELF-HARM, INIT
C2835428|T037|S22.078B|ICD10CM|OTHER FRACTURE OF T9-T10 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF T9-T10 VERTEBRA, INIT FOR OPN FX
C2835427|T037|S22.078A|ICD10CM|OTHER FRACTURE OF T9-T10 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF T9-T10 VERTEBRA, INIT FOR CLOS FX
C2877023|T037|T38.1X2S|ICD10CM|POISONING BY THYROID HORMONES AND SUBSTITUTES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY THYROID HORMONES AND SUB, SELF-HARM, SEQUELA
C2832299|T037|S06.359A|ICD10CM|TRAUMATIC HEMORRHAGE OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|TRAUM HEMOR LEFT CEREBRUM W LOC OF UNSP DURATION, INIT
C2832403|T037|S06.384A|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF BRAINSTEM WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|CONTUS/LAC/HEM BRAINSTEM W LOC OF 6 HOURS TO 24 HOURS, INIT
C2842142|T191|C50.929|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED SITE OF UNSPECIFIED MALE BREAST|MALIGNANT NEOPLASM OF UNSP SITE OF UNSPECIFIED MALE BREAST
C0238065|T047|K74.4|DMDICD10|SECONDARY BILIARY CIRRHOSIS|SEKUNDAERE BILIAERE ZIRRHOSE
C0023892|T047|K74.5|DMDICD10|BILIARY CIRRHOSIS, UNSPECIFIED|BILIAERE ZIRRHOSE, NICHT NAEHER BEZEICHNET
C0008312|T047|K74.3|DMDICD10|PRIMARY BILIARY CIRRHOSIS|PRIMAERE BILIAERE ZIRRHOSE
C2901804|T047|M86.139|ICD10CM|OTHER ACUTE OSTEOMYELITIS, UNSPECIFIED RADIUS AND ULNA|OTHER ACUTE OSTEOMYELITIS, UNSPECIFIED RADIUS AND ULNA
C2832405|T037|S06.384S|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF BRAINSTEM WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|CONTUS/LAC/HEM BRAINSTEM W LOC OF 6-24 HRS, SEQUELA
C2901803|T047|M86.132|ICD10CM|OTHER ACUTE OSTEOMYELITIS, LEFT RADIUS AND ULNA|OTHER ACUTE OSTEOMYELITIS, LEFT RADIUS AND ULNA
C2901802|T047|M86.131|ICD10CM|OTHER ACUTE OSTEOMYELITIS, RIGHT RADIUS AND ULNA|OTHER ACUTE OSTEOMYELITIS, RIGHT RADIUS AND ULNA
C2865552|T037|S88.119S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, UNSPECIFIED LOWER LEG, SEQUELA|COMPLETE TRAUM AMP AT LEV BETW KN & ANKL, UNSP LOW LEG, SQLA
C2878740|T037|T44.0X2S|ICD10CM|POISONING BY ANTICHOLINESTERASE AGENTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ANTICHOLINESTERASE AGENTS, SELF-HARM, SEQUELA
C2873898|T047|E08.319|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH UNSPECIFIED DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA|DIAB DUE TO UNDRL COND W UNSP DIAB RTNOP W/O MACULAR EDEMA
C3264212|T047|H40.1311|ICD10CM|PIGMENTARY GLAUCOMA, RIGHT EYE, MILD STAGE|PIGMENTARY GLAUCOMA, RIGHT EYE, MILD STAGE
C3264213|T047|H40.1312|ICD10CM|PIGMENTARY GLAUCOMA, RIGHT EYE, MODERATE STAGE|PIGMENTARY GLAUCOMA, RIGHT EYE, MODERATE STAGE
C3264214|T047|H40.1313|ICD10CM|PIGMENTARY GLAUCOMA, RIGHT EYE, SEVERE STAGE|PIGMENTARY GLAUCOMA, RIGHT EYE, SEVERE STAGE
C3264215|T047|H40.1314|ICD10CM|PIGMENTARY GLAUCOMA, RIGHT EYE, INDETERMINATE STAGE|PIGMENTARY GLAUCOMA, RIGHT EYE, INDETERMINATE STAGE
C2873897|T047|E08.311|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH UNSPECIFIED DIABETIC RETINOPATHY WITH MACULAR EDEMA|DIAB DUE TO UNDRL COND W UNSP DIABETIC RTNOP W MACULAR EDEMA
C2889283|T047|M05.551|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT HIP|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889284|T047|M05.552|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT HIP|RHEUMATOID POLYNEUROPATHY W RHEUMATOID ARTHRITIS OF LEFT HIP
C2842078|T191|C50.012|ICD10CM|MALIGNANT NEOPLASM OF NIPPLE AND AREOLA, LEFT FEMALE BREAST|MALIGNANT NEOPLASM OF NIPPLE AND AREOLA, LEFT FEMALE BREAST
C2878738|T037|T44.0X2A|ICD10CM|POISONING BY ANTICHOLINESTERASE AGENTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ANTICHOLINESTERASE AGENTS, SELF-HARM, INIT
C2865551|T037|S88.119D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, UNSPECIFIED LOWER LEG, SUBSEQUENT ENCOUNTER|COMPLETE TRAUM AMP AT LEV BETW KN & ANKL, UNSP LOW LEG, SUBS
C2837758|T037|S32.14XA|ICD10CM|TYPE 1 FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE 1 FRACTURE OF SACRUM, INIT ENCNTR FOR CLOSED FRACTURE
C2837759|T037|S32.14XB|ICD10CM|TYPE 1 FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE 1 FRACTURE OF SACRUM, INIT ENCNTR FOR OPEN FRACTURE
C0348484|T047|E71.19|ICD10CM|OTHER DISORDERS OF BRANCHED-CHAIN AMINO-ACID METABOLISM|OTHER DISORDERS OF BRANCHED-CHAIN AMINO-ACID METABOLISM
C2889295|T047|M05.59|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES|RHEUMATOID POLYNEUROPATHY W RHEUMATOID ARTHRITIS MULT SITE
C2896537|T046|M80.032A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, LEFT FOREARM, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, L FOREARM, INIT
C2889264|T047|M05.50|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP SITE
C2834040|T037|S14.153A|ICD10CM|OTHER INCOMPLETE LESION AT C3 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|OTH INCOMPLETE LESION AT C3, INIT
C2834041|T037|S14.153D|ICD10CM|OTHER INCOMPLETE LESION AT C3 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|OTH INCOMPLETE LESION AT C3, SUBS
C2889336|T047|M05.731|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT WRIST WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRITIS W RHEU FACTOR OF R WRIST W/O ORG/SYS INVOLV
C2889337|T047|M05.732|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT WRIST WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRITIS W RHEU FACTOR OF L WRIST W/O ORG/SYS INVOLV
C2889338|T047|M05.739|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED WRIST WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRIT W RHEU FACTOR OF UNSP WRIST W/O ORG/SYS INVOLV
C2834042|T037|S14.153S|ICD10CM|OTHER INCOMPLETE LESION AT C3 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|OTH INCOMPLETE LESION AT C3, SEQUELA
C2843303|T037|S48.119A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN UNSPECIFIED SHOULDER AND ELBOW, INITIAL ENCOUNTER|COMPLETE TRAUM AMP AT LEVEL BETW UNSP SHLDR AND ELBOW, INIT
C4269412|T037|S02.40FA|ICD10CM|ZYGOMATIC FRACTURE, LEFT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|ZYGOMATIC FRACTURE, LEFT SIDE, INIT
C2834011|T037|S14.145S|ICD10CM|BROWN-SEQUARD SYNDROME AT C5 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|BROWN-SEQUARD SYNDROME AT C5, SEQUELA
C2834009|T037|S14.145A|ICD10CM|BROWN-SEQUARD SYNDROME AT C5 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|BROWN-SEQUARD SYNDROME AT C5, INIT
C4269215|T033|R40.2444|ICD10CM|OTHER COMA, WITHOUT DOCUMENTED GLASGOW COMA SCALE SCORE, OR WITH PARTIAL SCORE REPORTED, 24 HOURS OR MORE AFTER HOSPITAL ADMISSION|OTHER COMA, WITHOUT GLASGOW, OR W/PART SCORE, 24+HRS
C4269214|T033|R40.2443|ICD10CM|OTHER COMA, WITHOUT DOCUMENTED GLASGOW COMA SCALE SCORE, OR WITH PARTIAL SCORE REPORTED, AT HOSPITAL ADMISSION|OTHER COMA, WITHOUT GLASGOW, OR W/PART SCORE, ADMIT
C4269213|T033|R40.2442|ICD10CM|OTHER COMA, WITHOUT DOCUMENTED GLASGOW COMA SCALE SCORE, OR WITH PARTIAL SCORE REPORTED, AT ARRIVAL TO EMERGENCY DEPARTMENT|OTHER COMA, WITHOUT DOCUMENTED GLASGOW, OR W/PART SCORE, EMR
C4269212|T033|R40.2441|ICD10CM|OTHER COMA, WITHOUT DOCUMENTED GLASGOW COMA SCALE SCORE, OR WITH PARTIAL SCORE REPORTED, IN THE FIELD [EMT OR AMBULANCE]|OTHER COMA, WITHOUT GLASGOW, OR W/PART SCORE, IN THE FIELD
C4269211|T033|R40.2440|ICD10CM|OTHER COMA, WITHOUT DOCUMENTED GLASGOW COMA SCALE SCORE, OR WITH PARTIAL SCORE REPORTED, UNSPECIFIED TIME|OTHER COMA, WITHOUT GLASGOW, OR W/PART SCORE, UNSP TIME
C0038663|T037|T14.91|ICD10CM|SUICIDE ATTEMPT|SUICIDE ATTEMPT
C2837459|T037|S32.002A|ICD10CM|UNSTABLE BURST FRACTURE OF UNSPECIFIED LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSTABLE BURST FRACTURE OF UNSP LUMBAR VERTEBRA, INIT
C4509256|T047|K56.50|ICD10CM|INTESTINAL ADHESIONS [BANDS], UNSPECIFIED AS TO PARTIAL VERSUS COMPLETE OBSTRUCTION|INTESTNL ADHESIONS, UNSP AS TO PARTIAL VERSUS COMPLETE OBST
C4509258|T047|K56.51|ICD10CM|INTESTINAL ADHESIONS [BANDS], WITH PARTIAL OBSTRUCTION|INTESTINAL ADHESIONS WITH INCOMPLETE OBSTRUCTION
C4509586|T047|K56.52|ICD10CM|INTESTINAL ADHESIONS [BANDS] WITH COMPLETE OBSTRUCTION|INTESTINAL ADHESIONS [BANDS] WITH COMPLETE OBSTRUCTION
C2891227|T037|T85.72XA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INSULIN PUMP, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INSULIN PUMP, INIT
C0694499|T047|I43|DMDICD10|CARDIOMYOPATHY IN DISEASES CLASSIFIED ELSEWHERE|KARDIOMYOPATHIE BEI ANDERENORTS KLASSIFIZIERTEN KRANKHEITEN
C2902121|T046|M87.376|ICD10CM|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED FOOT|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED FOOT
C2902122|T046|M87.377|ICD10CM|OTHER SECONDARY OSTEONECROSIS, RIGHT TOE(S)|OTHER SECONDARY OSTEONECROSIS, RIGHT TOE(S)
C2902119|T046|M87.374|ICD10CM|OTHER SECONDARY OSTEONECROSIS, RIGHT FOOT|OTHER SECONDARY OSTEONECROSIS, RIGHT FOOT
C2902120|T046|M87.375|ICD10CM|OTHER SECONDARY OSTEONECROSIS, LEFT FOOT|OTHER SECONDARY OSTEONECROSIS, LEFT FOOT
C2902117|T046|M87.372|ICD10CM|OTHER SECONDARY OSTEONECROSIS, LEFT ANKLE|OTHER SECONDARY OSTEONECROSIS, LEFT ANKLE
C2902118|T046|M87.373|ICD10CM|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED ANKLE|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED ANKLE
C2902116|T046|M87.371|ICD10CM|OTHER SECONDARY OSTEONECROSIS, RIGHT ANKLE|OTHER SECONDARY OSTEONECROSIS, RIGHT ANKLE
C0153377|T191|C05.2|DMDICD10|MALIGNANT NEOPLASM OF UVULA|BOESARTIGE NEUBILDUNG: UVULA
C2878408|T037|T43.222S|ICD10CM|POISONING BY SELECTIVE SEROTONIN REUPTAKE INHIBITORS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY SLCTV SEROTONIN REUPTAKE INHIBTR, SLF-HRM, SEQUELA
C2902123|T046|M87.378|ICD10CM|OTHER SECONDARY OSTEONECROSIS, LEFT TOE(S)|OTHER SECONDARY OSTEONECROSIS, LEFT TOE(S)
C2902124|T046|M87.379|ICD10CM|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED TOE(S)|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED TOE(S)
C4268043|T047|E10.3529|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, UNSPECIFIED EYE|TYPE 1 DIAB W PROLIF DIAB RTNOP WITH TRCTN DTCH MACULA, UNSP
C0837898|T047|M12.00|ICD10AM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], UNSPECIFIED SITE|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], MULTIPLE SITES
C2911426|T033|Z89.611|ICD10CM|ACQUIRED ABSENCE OF RIGHT LEG ABOVE KNEE|ACQUIRED ABSENCE OF RIGHT LEG ABOVE KNEE
C4268042|T047|E10.3523|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, BILATERAL|TYPE 1 DIAB W PROLIF DIAB RTNOP WITH TRCTN DTCH MACULA, BI
C4268041|T047|E10.3522|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, LEFT EYE|TYPE 1 DIAB W PROLIF DIAB RTNOP W TRCTN DTCH MACULA, L EYE
C4268040|T047|E10.3521|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, RIGHT EYE|TYPE 1 DIAB W PROLIF DIAB RTNOP W TRCTN DTCH MACULA, R EYE
C0837898|T047|M12.09|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], MULTIPLE SITES|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], MULTIPLE SITES
C3696796|T047|M12.08|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], OTHER SPECIFIED SITE|CHRONIC POSTRHEUMATIC ARTHROPATHY, OTHER SPECIFIED SITE
C2857890|T037|S72.335A|ICD10CM|NONDISPLACED OBLIQUE FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED OBLIQUE FRACTURE OF SHAFT OF LEFT FEMUR, INIT
C2860029|T037|S78.912S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT HIP AND THIGH, LEVEL UNSPECIFIED, SEQUELA|COMPLETE TRAUM AMP OF L HIP AND THIGH, LEVEL UNSP, SEQUELA
C2901046|T046|M84.464A|ICD10CM|PATHOLOGICAL FRACTURE, LEFT FIBULA, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, LEFT FIBULA, INIT ENCNTR FOR FRACTURE
C2859227|T037|S73.035A|ICD10CM|OTHER ANTERIOR DISLOCATION OF LEFT HIP, INITIAL ENCOUNTER|OTHER ANTERIOR DISLOCATION OF LEFT HIP, INITIAL ENCOUNTER
C2891205|T037|T85.691D|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTRAPERITONEAL DIALYSIS CATHETER, SUBSEQUENT ENCOUNTER|MECH COMPL OF INTRAPERITONEAL DIALYSIS CATHETER, SUBS ENCNTR
C2860028|T037|S78.912D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT HIP AND THIGH, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|COMPLETE TRAUM AMP OF LEFT HIP AND THIGH, LEVEL UNSP, SUBS
C2890662|T037|T84.191A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTERNAL FIXATION DEVICE OF LEFT HUMERUS, INITIAL ENCOUNTER|MECH COMPL OF INTERNAL FIXATION DEVICE OF LEFT HUMERUS, INIT
C2860027|T037|S78.912A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT HIP AND THIGH, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|COMPLETE TRAUM AMP OF LEFT HIP AND THIGH, LEVEL UNSP, INIT
C2865576|T037|S88.919A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED LOWER LEG, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMP OF UNSP LOWER LEG, LEVEL UNSP, INIT
C2890735|T037|T84.293A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTERNAL FIXATION DEVICE OF BONES OF FOOT AND TOES, INITIAL ENCOUNTER|MECH COMPL OF INT FIX OF BONES OF FOOT AND TOES, INIT
C2865577|T037|S88.919D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED LOWER LEG, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMP OF UNSP LOWER LEG, LEVEL UNSP, SUBS
C2901560|T046|M84.673A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, UNSPECIFIED ANKLE, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, UNSP ANKLE, INIT
C2865578|T037|S88.919S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED LOWER LEG, LEVEL UNSPECIFIED, SEQUELA|COMPLETE TRAUMATIC AMP OF UNSP LOW LEG, LEVEL UNSP, SEQUELA
C2877514|T037|T39.8X2S|ICD10CM|POISONING BY OTHER NONOPIOID ANALGESICS AND ANTIPYRETICS, NOT ELSEWHERE CLASSIFIED, INTENTIONAL SELF-HARM, SEQUELA|POISN BY OTH NONOPIO ANALGES/ANTIPYRET, NEC, SLF-HRM, SQLA
C4270250|T046|T83.112A|ICD10CM|BREAKDOWN (MECHANICAL) OF INDWELLING URETERAL STENT, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF INDWELLING URETERAL STENT, INIT
C2884762|T037|T58.12XA|ICD10CM|TOXIC EFFECT OF CARBON MONOXIDE FROM UTILITY GAS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CARB MONX FROM UTILITY GAS, SELF-HARM, INIT
C2860044|T037|S78.929A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED HIP AND THIGH, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|PARTIAL TRAUM AMP OF UNSP HIP AND THIGH, LEVEL UNSP, INIT
C2900954|T046|M84.442A|ICD10CM|PATHOLOGICAL FRACTURE, LEFT HAND, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, LEFT HAND, INIT ENCNTR FOR FRACTURE
C2900939|T046|M84.439A|ICD10CM|PATHOLOGICAL FRACTURE, UNSPECIFIED ULNA AND RADIUS, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, UNSP ULNA AND RADIUS, INIT FOR FX
C2888897|T047|M00.81|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, UNSPECIFIED SHOULDER|ARTHRITIS DUE TO OTHER BACTERIA, SHOULDER
C2900451|T047|A81.1|ICD10CM|SUBACUTE SCLEROSING PANENCEPHALITIS|VAN BOGAERT'S SCLEROSING LEUKOENCEPHALOPATHY
C0023524|T047|A81.2|DMDICD10|PROGRESSIVE MULTIFOCAL LEUKOENCEPHALOPATHY|PROGRESSIVE MULTIFOKALE LEUKENZEPHALOPATHIE
C2835758|T037|S24.101S|ICD10CM|UNSPECIFIED INJURY AT T1 LEVEL OF THORACIC SPINAL CORD, SEQUELA|UNSP INJURY AT T1 LEVEL OF THORACIC SPINAL CORD, SEQUELA
C2888896|T047|M00.812|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, LEFT SHOULDER|ARTHRITIS DUE TO OTHER BACTERIA, LEFT SHOULDER
C2888895|T047|M00.811|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, RIGHT SHOULDER|ARTHRITIS DUE TO OTHER BACTERIA, RIGHT SHOULDER
C0851226|T047|A81|ICD10CM|ATYPICAL VIRUS INFECTION OF CENTRAL NERVOUS SYSTEM, UNSPECIFIED|ATYPICAL VIRUS INFECTIONS OF CENTRAL NERVOUS SYSTEM
C2882926|T047|I70.619|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, UNSPECIFIED EXTREMITY|ATHSCL NONBIOL BYPASS OF EXTRM W INTRMT CLAUD, UNSP EXTRM
C2882925|T047|I70.618|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, OTHER EXTREMITY|ATHSCL NONBIOL BYPASS OF THE EXTRM W INTRMT CLAUD, OTH EXTRM
C2882924|T047|I70.613|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, BILATERAL LEGS|ATHSCL NONBIOL BYPASS OF THE EXTRM W INTRMT CLAUD, BI LEGS
C2882923|T047|I70.612|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, LEFT LEG|ATHSCL NONBIOL BYPASS OF THE EXTRM W INTRMT CLAUD, LEFT LEG
C2882922|T047|I70.611|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH INTERMITTENT CLAUDICATION, RIGHT LEG|ATHSCL NONBIOL BYPASS OF THE EXTRM W INTRMT CLAUD, RIGHT LEG
C2835855|T037|S24.154S|ICD10CM|OTHER INCOMPLETE LESION AT T11-T12 LEVEL OF THORACIC SPINAL CORD, SEQUELA|OTH INCOMPLETE LESION AT T11-T12, SEQUELA
C2854052|T191|C85.89|ICD10CM|OTHER SPECIFIED TYPES OF NON-HODGKIN LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES|OTH TYPES OF NON-HODG LYMPH, EXTRNOD AND SOLID ORGAN SITES
C2854051|T191|C85.88|ICD10CM|OTHER SPECIFIED TYPES OF NON-HODGKIN LYMPHOMA, LYMPH NODES OF MULTIPLE SITES|OTH TYPES OF NON-HODGKIN LYMPHOMA, LYMPH NODES MULT SITE
C2901140|T046|M84.511A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, RIGHT SHOULDER, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, R SHOULDER, INIT
C2854046|T191|C85.83|ICD10CM|OTHER SPECIFIED TYPES OF NON-HODGKIN LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES|OTH TYPES OF NON-HODGKIN LYMPHOMA, INTRA-ABD LYMPH NODES
C2854045|T191|C85.82|ICD10CM|OTHER SPECIFIED TYPES OF NON-HODGKIN LYMPHOMA, INTRATHORACIC LYMPH NODES|OTH TYPES OF NON-HODGKIN LYMPHOMA, INTRATHORACIC LYMPH NODES
C2854044|T191|C85.81|ICD10CM|OTHER SPECIFIED TYPES OF NON-HODGKIN LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK|OTH TYPES OF NON-HODG LYMPH, NODES OF HEAD, FACE, AND NECK
C2854043|T191|C85.80|ICD10CM|OTHER SPECIFIED TYPES OF NON-HODGKIN LYMPHOMA, UNSPECIFIED SITE|OTH TYPES OF NON-HODGKIN LYMPHOMA, UNSPECIFIED SITE
C2854050|T191|C85.87|ICD10CM|OTHER SPECIFIED TYPES OF NON-HODGKIN LYMPHOMA, SPLEEN|OTHER SPECIFIED TYPES OF NON-HODGKIN LYMPHOMA, SPLEEN
C2854049|T191|C85.86|ICD10CM|OTHER SPECIFIED TYPES OF NON-HODGKIN LYMPHOMA, INTRAPELVIC LYMPH NODES|OTH TYPES OF NON-HODGKIN LYMPHOMA, INTRAPELVIC LYMPH NODES
C2854048|T191|C85.85|ICD10CM|OTHER SPECIFIED TYPES OF NON-HODGKIN LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|OTH TYPES OF NON-HODG LYMPH, NODES OF ING RGN AND LOWER LIMB
C2854047|T191|C85.84|ICD10CM|OTHER SPECIFIED TYPES OF NON-HODGKIN LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB|OTH TYPES OF NON-HODG LYMPH, NODES OF AXILLA AND UPPER LIMB
C0345904|T191|C22.9|DMDICD10|MALIGNANT NEOPLASM OF LIVER, NOT SPECIFIED AS PRIMARY OR SECONDARY|BOESARTIGE NEUBILDUNG: LEBER, NICHT NAEHER BEZEICHNET
C2837938|T191|C22.8|ICD10CM|MALIGNANT NEOPLASM OF LIVER, PRIMARY, UNSPECIFIED AS TO TYPE|MALIGNANT NEOPLASM OF LIVER, PRIMARY, UNSPECIFIED AS TO TYPE
C0348339|T191|C22.4|DMDICD10|OTHER SARCOMAS OF LIVER|SONSTIGE SARKOME DER LEBER
C0348340|T191|C22.7|DMDICD10|OTHER SPECIFIED CARCINOMAS OF LIVER|SONSTIGE NAEHER BEZEICHNETE KARZINOME DER LEBER
C2857634|T037|S72.25XC|ICD10CM|NONDISPLACED SUBTROCHANTERIC FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP SUBTROCHNT FX L FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C0345905|T191|C22.1|DMDICD10|INTRAHEPATIC BILE DUCT CARCINOMA|INTRAHEPATISCHES GALLENGANGSKARZINOM
C2239176|T191|C22.0|DMDICD10|LIVER CELL CARCINOMA|LEBERZELLKARZINOM
C0345907|T191|C22.3|DMDICD10|ANGIOSARCOMA OF LIVER|ANGIOSARKOM DER LEBER
C0206624|T191|C22.2|DMDICD10|HEPATOBLASTOMA|HEPATOBLASTOM
C2901883|T047|M86.459|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, UNSPECIFIED FEMUR|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, UNSPECIFIED FEMUR
C2832080|T037|S06.306S|ICD10CM|UNSPECIFIED FOCAL TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|UNSP FOCAL TBI W LOC >24 HR W/O RET CONSC W SURV, SEQUELA
C2890778|T037|T84.418A|ICD10CM|BREAKDOWN (MECHANICAL) OF OTHER INTERNAL ORTHOPEDIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|BRKDWN INTERNAL ORTH DEVICES, IMPLANTS AND GRAFTS, INIT
C2901881|T047|M86.451|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, RIGHT FEMUR|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, RIGHT FEMUR
C2901882|T047|M86.452|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, LEFT FEMUR|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, LEFT FEMUR
C2832078|T037|S06.306A|ICD10CM|UNSPECIFIED FOCAL TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|UNSP FOCAL TBI W LOC >24 HR W/O RET CONSC W SURV, INIT
C2879257|T037|T45.622A|ICD10CM|POISONING BY HEMOSTATIC DRUG, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY HEMOSTATIC DRUG, INTENTIONAL SELF-HARM, INIT
C2858968|T037|S72.479A|ICD10CM|TORUS FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TORUS FRACTURE OF LOWER END OF UNSP FEMUR, INIT FOR CLOS FX
C2855838|T037|S68.011S|ICD10CM|COMPLETE TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF RIGHT THUMB, SEQUELA|COMPLETE TRAUMATIC MCP AMPUTATION OF RIGHT THUMB, SEQUELA
C2869824|T037|S98.142A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF ONE LEFT LESSER TOE, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF ONE LEFT LESSER TOE, INIT
C2869825|T037|S98.142D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF ONE LEFT LESSER TOE, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF ONE LEFT LESSER TOE, SUBS
C2833859|T037|S14.104D|ICD10CM|UNSPECIFIED INJURY AT C4 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY AT C4 LEVEL OF CERVICAL SPINAL CORD, SUBS ENCNTR
C2869826|T037|S98.142S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF ONE LEFT LESSER TOE, SEQUELA|PARTIAL TRAUMATIC AMPUTATION OF ONE LEFT LESSER TOE, SEQUELA
C2349509|T047||ICD10CM|CORONARY ATHEROSCLEROSIS DUE TO LIPID RICH PLAQUE
C1955780|T047|I25.82|ICD10CM|CHRONIC TOTAL OCCLUSION OF CORONARY ARTERY|TOTAL OCCLUSION OF CORONARY ARTERY
C2842154|T191|C57.20|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED ROUND LIGAMENT|MALIGNANT NEOPLASM OF UNSPECIFIED ROUND LIGAMENT
C2842155|T191|C57.21|ICD10CM|MALIGNANT NEOPLASM OF RIGHT ROUND LIGAMENT|MALIGNANT NEOPLASM OF RIGHT ROUND LIGAMENT
C2842156|T191|C57.22|ICD10CM|MALIGNANT NEOPLASM OF LEFT ROUND LIGAMENT|MALIGNANT NEOPLASM OF LEFT ROUND LIGAMENT
C3161193|T047|I25.84|ICD10CM|CORONARY ATHEROSCLEROSIS DUE TO CALCIFIED CORONARY LESION|CORONARY ATHEROSCLEROSIS DUE TO SEVERELY CALCIFIED CORONARY LESION
C0155669|T047|I25.8|ICD10CM|OTHER FORMS OF CHRONIC ISCHEMIC HEART DISEASE|OTHER FORMS OF CHRONIC ISCHEMIC HEART DISEASE
C2833858|T037|S14.104A|ICD10CM|UNSPECIFIED INJURY AT C4 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY AT C4 LEVEL OF CERVICAL SPINAL CORD, INIT ENCNTR
C2890898|T037|T84.81XA|ICD10CM|EMBOLISM DUE TO INTERNAL ORTHOPEDIC PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|EMBOLISM DUE TO INTERNAL ORTHOPEDIC PROSTH DEV/GRFT, INIT
C2857274|T037|S72.122A|ICD10CM|DISPLACED FRACTURE OF LESSER TROCHANTER OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF LESSER TROCHANTER OF LEFT FEMUR, INIT FOR CLOS FX
C2857275|T037|S72.122B|ICD10CM|DISPLACED FRACTURE OF LESSER TROCHANTER OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF LESS TROCHANTER OF L FEMR, 7THB
C2857276|T037|S72.122C|ICD10CM|DISPLACED FRACTURE OF LESSER TROCHANTER OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF LESS TROCHANTER OF L FEMR, 7THC
C2874904|T048|F31.76|ICD10CM|BIPOLAR DISORDER, IN FULL REMISSION, MOST RECENT EPISODE DEPRESSED|BIPOLAR DISORDER, IN FULL REMIS, MOST RECENT EPISODE DEPRESS
C2874905|T048|F31.77|ICD10CM|BIPOLAR DISORDER, IN PARTIAL REMISSION, MOST RECENT EPISODE MIXED|BIPOLAR DISORD, IN PARTIAL REMIS, MOST RECENT EPISODE MIXED
C2874902|T048|F31.74|ICD10CM|BIPOLAR DISORDER, IN FULL REMISSION, MOST RECENT EPISODE MANIC|BIPOLAR DISORDER, IN FULL REMIS, MOST RECENT EPISODE MANIC
C2874903|T048|F31.75|ICD10CM|BIPOLAR DISORDER, IN PARTIAL REMISSION, MOST RECENT EPISODE DEPRESSED|BIPOLAR DISORD, IN PARTIAL REMIS, MOST RECENT EPSD DEPRESS
C2874900|T048|F31.72|ICD10CM|BIPOLAR DISORDER, IN FULL REMISSION, MOST RECENT EPISODE HYPOMANIC|BIPOLAR DISORD, IN FULL REMIS, MOST RECENT EPISODE HYPOMANIC
C2874901|T048|F31.73|ICD10CM|BIPOLAR DISORDER, IN PARTIAL REMISSION, MOST RECENT EPISODE MANIC|BIPOLAR DISORD, IN PARTIAL REMIS, MOST RECENT EPISODE MANIC
C2874898|T048|F31.70|ICD10CM|BIPOLAR DISORDER, CURRENTLY IN REMISSION, MOST RECENT EPISODE UNSPECIFIED|BIPOLAR DISORD, CURRENTLY IN REMIS, MOST RECENT EPISODE UNSP
C2874899|T048|F31.71|ICD10CM|BIPOLAR DISORDER, IN PARTIAL REMISSION, MOST RECENT EPISODE HYPOMANIC|BIPOLAR DISORD, IN PARTIAL REMIS, MOST RECENT EPSD HYPOMANIC
C2874906|T048|F31.78|ICD10CM|BIPOLAR DISORDER, IN FULL REMISSION, MOST RECENT EPISODE MIXED|BIPOLAR DISORDER, IN FULL REMIS, MOST RECENT EPISODE MIXED
C0694525|T047|N08|DMDICD10|GLOMERULAR DISORDERS IN DISEASES CLASSIFIED ELSEWHERE|GLOMERULAERE KRANKHEITEN BEI ANDERENORTS KLASSIFIZIERTEN KRANKHEITEN
C2521617|T060|C23|ICD10PCS|MALIGNANT NEOPLASM OF GALLBLADDER|NUCLEAR MEDICINE, HEART, PET IMAG
C0949022|T191|C20|DMDICD10|MALIGNANT NEOPLASM OF RECTUM|BOESARTIGE NEUBILDUNG DES REKTUMS
C2882292|T047|I60.02|ICD10CM|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM LEFT CAROTID SIPHON AND BIFURCATION|NTRM SUBARACH HEMORRHAGE FROM LEFT CAROTID SIPHON AND BIFURC
C2882290|T047|I60.00|ICD10CM|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM UNSPECIFIED CAROTID SIPHON AND BIFURCATION|NTRM SUBARACH HEMORRHAGE FROM UNSP CAROTID SIPHON AND BIFURC
C2882291|T047|I60.01|ICD10CM|NONTRAUMATIC SUBARACHNOID HEMORRHAGE FROM RIGHT CAROTID SIPHON AND BIFURCATION|NTRM SUBARACH HEMOR FROM RIGHT CAROTID SIPHON AND BIFURC
C2832487|T037|S06.5X4S|ICD10CM|TRAUMATIC SUBDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|TRAUM SUBDR HEM W LOC OF 6 HOURS TO 24 HOURS, SEQUELA
C2890922|T037|T84.89XA|ICD10CM|OTHER SPECIFIED COMPLICATION OF INTERNAL ORTHOPEDIC PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|OTH COMP OF INTERNAL ORTHOPEDIC PROSTH DEV/GRFT, INIT
C2874435|T048|F11.19|ICD10CM|OPIOID ABUSE WITH UNSPECIFIED OPIOID-INDUCED DISORDER|OPIOID ABUSE WITH UNSPECIFIED OPIOID-INDUCED DISORDER
C4268215|T048|F11.14|ICD10CM|OPIOID ABUSE WITH OPIOID-INDUCED MOOD DISORDER|OPIOID USE DISORDER, MILD, WITH OPIOID-INDUCED DEPRESSIVE DISORDER
C2832485|T037|S06.5X4A|ICD10CM|TRAUMATIC SUBDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|TRAUM SUBDR HEM W LOC OF 6 HOURS TO 24 HOURS, INIT
C2832240|T037|S06.345A|ICD10CM|TRAUMATIC HEMORRHAGE OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, INITIAL ENCOUNTER|TRAUM HEMOR R CEREB W LOC >24 HR W RET CONSC LEV, INIT
C2838647|T037|S34.112S|ICD10CM|COMPLETE LESION OF L2 LEVEL OF LUMBAR SPINAL CORD, SEQUELA|COMPLETE LESION OF L2 LEVEL OF LUMBAR SPINAL CORD, SEQUELA
C2859252|T037|S73.045A|ICD10CM|CENTRAL DISLOCATION OF LEFT HIP, INITIAL ENCOUNTER|CENTRAL DISLOCATION OF LEFT HIP, INITIAL ENCOUNTER
C2895339|T037|M48.57XA|ICD10CM|COLLAPSED VERTEBRA, NOT ELSEWHERE CLASSIFIED, LUMBOSACRAL REGION, INITIAL ENCOUNTER FOR FRACTURE|COLLAPSED VERTEBRA, NEC, LUMBOSACRAL REGION, INIT
C2901919|T047|M86.631|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, RIGHT RADIUS AND ULNA|OTHER CHRONIC OSTEOMYELITIS, RIGHT RADIUS AND ULNA
C2901920|T047|M86.632|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, LEFT RADIUS AND ULNA|OTHER CHRONIC OSTEOMYELITIS, LEFT RADIUS AND ULNA
C2902081|T046|M87.31|ICD10CM|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED SHOULDER|OTHER SECONDARY OSTEONECROSIS, SHOULDER
C2833860|T037|S14.104S|ICD10CM|UNSPECIFIED INJURY AT C4 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|UNSP INJURY AT C4 LEVEL OF CERVICAL SPINAL CORD, SEQUELA
C2901921|T047|M86.639|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, UNSPECIFIED RADIUS AND ULNA|OTHER CHRONIC OSTEOMYELITIS, UNSPECIFIED RADIUS AND ULNA
C2890521|T037|T84.058A|ICD10CM|PERIPROSTHETIC OSTEOLYSIS OF OTHER INTERNAL PROSTHETIC JOINT, INITIAL ENCOUNTER|PERIPROSTHETIC OSTEOLYSIS OF INTERNAL PROSTHETIC JOINT, INIT
C2882277|T047|I50.9|ICD10CM|HEART FAILURE, UNSPECIFIED|CARDIAC, HEART OR MYOCARDIAL FAILURE NOS
C2889569|T047|M08.27|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, UNSPECIFIED ANKLE AND FOOT|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, ANKLE AND FOOT
C2857429|T037|S72.135B|ICD10CM|NONDISPLACED APOPHYSEAL FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP APOPHYSEAL FX LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C4509222|T047|I50.1|ICD10CM|LEFT VENTRICULAR FAILURE, UNSPECIFIED|LEFT VENTRICULAR FAILURE, UNSPECIFIED
C2889571|T047|M08.272|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, LEFT ANKLE AND FOOT|JUVENILE RHEUMATOID ARTHRITIS W SYSTEMIC ONSET, LEFT ANK/FT
C2889570|T047|M08.271|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, RIGHT ANKLE AND FOOT|JUVENILE RHEUMATOID ARTHRITIS W SYSTEMIC ONSET, RIGHT ANK/FT
C2888879|T047|M00.251|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, RIGHT HIP|OTHER STREPTOCOCCAL ARTHRITIS, RIGHT HIP
C2888880|T047|M00.252|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, LEFT HIP|OTHER STREPTOCOCCAL ARTHRITIS, LEFT HIP
C2832551|T037|S06.810S|ICD10CM|INJURY OF RIGHT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|INJURY OF R INT CAROTID, INTCR W/O LOC, SEQUELA
C2888881|T047|M00.259|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, UNSPECIFIED HIP|OTHER STREPTOCOCCAL ARTHRITIS, UNSPECIFIED HIP
C2857430|T037|S72.135C|ICD10CM|NONDISPLACED APOPHYSEAL FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP APOPHYSEAL FX L FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2832549|T037|S06.810A|ICD10CM|INJURY OF RIGHT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|INJURY OF R INT CAROTID, INTCR W/O LOC, INIT
C2886732|T037|T79.4XXA|ICD10CM|TRAUMATIC SHOCK, INITIAL ENCOUNTER|TRAUMATIC SHOCK, INITIAL ENCOUNTER
C2889528|T047|M08.01|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED SHOULDER|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, SHOULDER
C2889527|T047|M08.012|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, LEFT SHOULDER|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, LEFT SHOULDER
C2887264|T047|I85.10|ICD10CM|SECONDARY ESOPHAGEAL VARICES WITHOUT BLEEDING|SECONDARY ESOPHAGEAL VARICES WITHOUT BLEEDING
C2887265|T020|I85.11|ICD10CM|SECONDARY ESOPHAGEAL VARICES WITH BLEEDING|SECONDARY ESOPHAGEAL VARICES WITH BLEEDING
C2837596|T037|S32.041A|ICD10CM|STABLE BURST FRACTURE OF FOURTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|STABLE BURST FRACTURE OF FOURTH LUMBAR VERTEBRA, INIT
C2837597|T037|S32.041B|ICD10CM|STABLE BURST FRACTURE OF FOURTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|STABLE BURST FX FOURTH LUM VERTEBRA, INIT FOR OPN FX
C4509468|T037|T14.91XD|ICD10CM|SUICIDE ATTEMPT, SUBSEQUENT ENCOUNTER|SUICIDE ATTEMPT, SUBSEQUENT ENCOUNTER
C2832445|T037|S06.4X4A|ICD10CM|EPIDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|EPIDURAL HEMORRHAGE W LOC OF 6 HOURS TO 24 HOURS, INIT
C4509467|T037|T14.91XA|ICD10CM|SUICIDE ATTEMPT, INITIAL ENCOUNTER|SUICIDE ATTEMPT, INITIAL ENCOUNTER
C2886330|T037|T71.112A|ICD10CM|ASPHYXIATION DUE TO SMOTHERING UNDER PILLOW, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|ASPHYXIATION DUE TO SMOTHERING UNDER PILLOW, SELF-HARM, INIT
C2832447|T037|S06.4X4S|ICD10CM|EPIDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|EPIDURAL HEMORRHAGE W LOC OF 6 HOURS TO 24 HOURS, SEQUELA
C2890280|T037|T83.190A|ICD10CM|OTHER MECHANICAL COMPLICATION OF URINARY ELECTRONIC STIMULATOR DEVICE, INITIAL ENCOUNTER|MECH COMPL OF URINARY ELECTRONIC STIMULATOR DEVICE, INIT
C2860237|T037|S79.192A|ICD10CM|OTHER PHYSEAL FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH PHYSEAL FRACTURE OF LOWER END OF LEFT FEMUR, INIT
C2886332|T037|T71.112S|ICD10CM|ASPHYXIATION DUE TO SMOTHERING UNDER PILLOW, INTENTIONAL SELF-HARM, SEQUELA|ASPHYX DUE TO SMOTHERING UNDER PILLOW, SELF-HARM, SEQUELA
C3469322|T047|M05.059|ICD10CM|FELTY'S SYNDROME, UNSPECIFIED HIP|FELTY'S SYNDROME, UNSPECIFIED HIP
C2888930|T047|M01.X12|ICD10CM|DIRECT INFECTION OF LEFT SHOULDER IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIRECT INFCT OF L SHLDR IN INFEC/PARASTC DIS CLASSD ELSWHR
C2888931|T047|M01.X19|ICD10CM|DIRECT INFECTION OF UNSPECIFIED SHOULDER IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIR INFCT OF UNSP SHLDR IN INFEC/PARASTC DIS CLASSD ELSWHR
C2889123|T047|M05.052|ICD10CM|FELTY'S SYNDROME, LEFT HIP|FELTY'S SYNDROME, LEFT HIP
C2860003|T037|S78.112S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN LEFT HIP AND KNEE, SEQUELA|COMPLETE TRAUM AMP AT LEVEL BETW LEFT HIP AND KNEE, SEQUELA
C2833302|T037|S12.190B|ICD10CM|OTHER DISPLACED FRACTURE OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH DISP FX OF SECOND CERVICAL VERTEBRA, INIT FOR OPN FX
C2879519|T037|T46.5X2S|ICD10CM|POISONING BY OTHER ANTIHYPERTENSIVE DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH ANTIHYPERTENSIVE DRUGS, SELF-HARM, SEQUELA
C2860002|T037|S78.112D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN LEFT HIP AND KNEE, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMP AT LEVEL BETW LEFT HIP AND KNEE, SUBS
C2860001|T037|S78.112A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN LEFT HIP AND KNEE, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMP AT LEVEL BETW LEFT HIP AND KNEE, INIT
C2832142|T037|S06.321S|ICD10CM|CONTUSION AND LACERATION OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|CONTUS/LAC L CEREB W LOC OF 30 MINUTES OR LESS, SEQUELA
C4270311|T046|T83.510A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO CYSTOSTOMY CATHETER, INITIAL ENCOUNTER|I/I REACT D/T CYSTOSTOMY CATHETER, INITIAL ENCOUNTER
C2889385|T047|M05|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR, UNSPECIFIED|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR
C4269503|T037|S02.640A|ICD10CM|FRACTURE OF RAMUS OF MANDIBLE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF RAMUS OF MANDIBLE, UNSPECIFIED SIDE, INIT
C4268019|T047|E10.3311|ICD10CM|TYPE 1 DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|TYPE 1 DIAB WITH MOD NONP RTNOP WITH MACULAR EDEMA, R EYE
C4268020|T047|E10.3312|ICD10CM|TYPE 1 DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|TYPE 1 DIAB WITH MOD NONP RTNOP WITH MACULAR EDEMA, L EYE
C4268021|T047|E10.3313|ICD10CM|TYPE 1 DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|TYPE 1 DIAB WITH MODERATE NONP RTNOP WITH MACULAR EDEMA, BI
C4269504|T037|S02.640B|ICD10CM|FRACTURE OF RAMUS OF MANDIBLE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF RAMUS OF MANDIBLE, UNSPECIFIED SIDE, 7THB
C2832140|T037|S06.321A|ICD10CM|CONTUSION AND LACERATION OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|CONTUS/LAC LEFT CEREBRUM W LOC OF 30 MINUTES OR LESS, INIT
C2902007|T046|M87.145|ICD10CM|OSTEONECROSIS DUE TO DRUGS, LEFT FINGER(S)|OSTEONECROSIS DUE TO DRUGS, LEFT FINGER(S)
C4268022|T047|E10.3319|ICD10CM|TYPE 1 DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|TYPE 1 DIAB WITH MOD NONP RTNOP WITH MACULAR EDEMA, UNSP
C2902008|T046|M87.146|ICD10CM|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED FINGER(S)|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED FINGER(S)
C2902003|T046|M87.141|ICD10CM|OSTEONECROSIS DUE TO DRUGS, RIGHT HAND|OSTEONECROSIS DUE TO DRUGS, RIGHT HAND
C2902005|T046|M87.143|ICD10CM|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED HAND|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED HAND
C2902004|T046|M87.142|ICD10CM|OSTEONECROSIS DUE TO DRUGS, LEFT HAND|OSTEONECROSIS DUE TO DRUGS, LEFT HAND
C2865591|T037|S88.929S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED LOWER LEG, LEVEL UNSPECIFIED, SEQUELA|PARTIAL TRAUMATIC AMP OF UNSP LOWER LEG, LEVEL UNSP, SEQUELA
C2856692|T037|S72.031C|ICD10CM|DISPLACED MIDCERVICAL FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL MIDCERVICAL FX R FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C0341102|T047|K21.9|DMDICD10|GASTRO-ESOPHAGEAL REFLUX DISEASE WITHOUT ESOPHAGITIS|GASTROOESOPHAGEALE REFLUXKRANKHEIT OHNE OESOPHAGITIS
C2856690|T037|S72.031A|ICD10CM|DISPLACED MIDCERVICAL FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED MIDCERVICAL FRACTURE OF RIGHT FEMUR, INIT
C2902125|T046|M87.80|ICD10CM|OTHER OSTEONECROSIS, UNSPECIFIED BONE|OTHER OSTEONECROSIS, UNSPECIFIED BONE
C0677659|T047|K21.0|DMDICD10|GASTRO-ESOPHAGEAL REFLUX DISEASE WITH ESOPHAGITIS|GASTROOESOPHAGEALE REFLUXKRANKHEIT MIT OESOPHAGITIS
C1384514|T047||ICD10CM|CONN'S SYNDROME
C1260386|T047|E26.02|ICD10CM|GLUCOCORTICOID-REMEDIABLE ALDOSTERONISM|GLUCOCORTICOID-REMEDIABLE ALDOSTERONISM
C0840057|T046|M87.88|ICD10AM|OTHER OSTEONECROSIS, OTHER SITE|OTHER OSTEONECROSIS, OTHER SITE
C4269580|T037|S02.82XA|ICD10CM|FRACTURE OF OTHER SPECIFIED SKULL AND FACIAL BONES, LEFT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF OTH SKULL AND FACIAL BONES, LEFT SIDE, INIT
C4269581|T037|S02.82XB|ICD10CM|FRACTURE OF OTHER SPECIFIED SKULL AND FACIAL BONES, LEFT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF OTH SKULL AND FACIAL BONES, LEFT SIDE, 7THB
C2901132|T046|M84.50XA|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, UNSPECIFIED SITE, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, UNSP SITE, INIT
C2902854|T047|N00.8|ICD10CM|ACUTE NEPHRITIC SYNDROME WITH OTHER MORPHOLOGIC CHANGES|ACUTE NEPHRITIC SYNDROME WITH OTHER MORPHOLOGIC CHANGES
C2889112|T047|M05.021|ICD10CM|FELTY'S SYNDROME, RIGHT ELBOW|FELTY'S SYNDROME, RIGHT ELBOW
C2902851|T047|N00.6|ICD10CM|ACUTE NEPHRITIC SYNDROME WITH DENSE DEPOSIT DISEASE|ACUTE NEPHRITIC SYNDROME WITH MEMBRANOPROLIFERATIVE GLOMERULONEPHRITIS, TYPE 2
C2902852|T047|N00.7|ICD10CM|ACUTE NEPHRITIC SYNDROME WITH DIFFUSE CRESCENTIC GLOMERULONEPHRITIS|ACUTE NEPHRITIC SYNDROME WITH EXTRACAPILLARY GLOMERULONEPHRITIS
C0451741|T047|N00.4|DMDICD10|ACUTE NEPHRITIC SYNDROME WITH DIFFUSE ENDOCAPILLARY PROLIFERATIVE GLOMERULONEPHRITIS|AKUTES NEPHRITISCHES SYNDROM: DIFFUSE ENDOKAPILLAER-PROLIFERATIVE GLOMERULONEPHRITIS
C2902850|T047|N00.5|ICD10CM|ACUTE NEPHRITIC SYNDROME WITH DIFFUSE MESANGIOCAPILLARY GLOMERULONEPHRITIS|ACUTE NEPHRITIC SYNDROME WITH MEMBRANOPROLIFERATIVE GLOMERULONEPHRITIS, TYPES 1 AND 3, OR NOS
C0451739|T047|N00.2|DMDICD10|ACUTE NEPHRITIC SYNDROME WITH DIFFUSE MEMBRANOUS GLOMERULONEPHRITIS|AKUTES NEPHRITISCHES SYNDROM: DIFFUSE MEMBRANOESE GLOMERULONEPHRITIS
C0451740|T047|N00.3|DMDICD10|ACUTE NEPHRITIC SYNDROME WITH DIFFUSE MESANGIAL PROLIFERATIVE GLOMERULONEPHRITIS|AKUTES NEPHRITISCHES SYNDROM: DIFFUSE MESANGIOPROLIFERATIVE GLOMERULONEPHRITIS
C2902846|T047|N00.0|ICD10CM|ACUTE NEPHRITIC SYNDROME WITH MINOR GLOMERULAR ABNORMALITY|ACUTE NEPHRITIC SYNDROME WITH MINIMAL CHANGE LESION
C2902849|T047|N00.1|ICD10CM|ACUTE NEPHRITIC SYNDROME WITH FOCAL AND SEGMENTAL GLOMERULAR LESIONS|ACUTE NEPHRITIC SYNDROME WITH FOCAL GLOMERULONEPHRITIS
C2838136|T037|S32.441A|ICD10CM|DISPLACED FRACTURE OF POSTERIOR COLUMN [ILIOISCHIAL] OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF POSTERIOR COLUMN OF RIGHT ACETABULUM, INIT
C2838137|T037|S32.441B|ICD10CM|DISPLACED FRACTURE OF POSTERIOR COLUMN [ILIOISCHIAL] OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISP FX OF POSTERIOR COLUMN OF RIGHT ACETAB, INIT FOR OPN FX
C4268067|T047|E10.37X9|ICD10CM|TYPE 1 DIABETES MELLITUS WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, UNSPECIFIED EYE|TYPE 1 DIAB WITH DIAB MCLR EDEMA, RESOLVED FOL TRTMT, UNSP
C4268066|T047|E10.37X3|ICD10CM|TYPE 1 DIABETES MELLITUS WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, BILATERAL|TYPE 1 DIAB WITH DIAB MACULAR EDEMA, RESOLVED FOL TRTMT, BI
C4268065|T047|E10.37X2|ICD10CM|TYPE 1 DIABETES MELLITUS WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, LEFT EYE|TYPE 1 DIAB WITH DIAB MCLR EDEMA, RESOLVED FOL TRTMT, L EYE
C4268064|T047|E10.37X1|ICD10CM|TYPE 1 DIABETES MELLITUS WITH DIABETIC MACULAR EDEMA, RESOLVED FOLLOWING TREATMENT, RIGHT EYE|TYPE 1 DIAB WITH DIAB MCLR EDEMA, RESOLVED FOL TRTMT, R EYE
C4509265|T047|K56.691|ICD10CM|OTHER COMPLETE INTESTINAL OBSTRUCTION|OTHER COMPLETE INTESTINAL OBSTRUCTION
C4509264|T047|K56.690|ICD10CM|OTHER PARTIAL INTESTINAL OBSTRUCTION|OTHER INCOMPLETE INTESTINAL OBSTRUCTION
C2977855|T037|S32.509A|ICD10CM|UNSPECIFIED FRACTURE OF UNSPECIFIED PUBIS, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF UNSP PUBIS, INIT ENCNTR FOR CLOSED FRACTURE
C4509267|T047|K56.699|ICD10CM|OTHER INTESTINAL OBSTRUCTION UNSPECIFIED AS TO PARTIAL VERSUS COMPLETE OBSTRUCTION|OTHER INTESTINAL OBSTRUCTION, NEC
C2856019|T037|S68.614S|ICD10CM|COMPLETE TRAUMATIC TRANSPHALANGEAL AMPUTATION OF RIGHT RING FINGER, SEQUELA|COMPLETE TRAUMATIC TRNSPHAL AMP OF R RNG FNGR, SEQUELA
C2877537|T037|T39.92XA|ICD10CM|POISONING BY UNSPECIFIED NONOPIOID ANALGESIC, ANTIPYRETIC AND ANTIRHEUMATIC, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY UNSP NONOPI ANALGS/ANTIPYR/ANTIRHEU, SLF-HRM, INIT
C2884802|T037|T58.8X2S|ICD10CM|TOXIC EFFECT OF CARBON MONOXIDE FROM OTHER SOURCE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CARB MONX FROM OTH SOURCE, SLF-HRM, SEQUELA
C2837949|T191|C34.02|ICD10CM|MALIGNANT NEOPLASM OF LEFT MAIN BRONCHUS|MALIGNANT NEOPLASM OF LEFT MAIN BRONCHUS
C2845906|T191|C69.21|ICD10CM|MALIGNANT NEOPLASM OF RIGHT RETINA|MALIGNANT NEOPLASM OF RIGHT RETINA
C2858645|T037|S72.441B|ICD10CM|DISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF LOW EPIPHY (SEPARATION) OF R FEMR, 7THB
C2858646|T037|S72.441C|ICD10CM|DISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF LOW EPIPHY (SEPARATION) OF R FEMR, 7THC
C2877539|T037|T39.92XS|ICD10CM|POISONING BY UNSPECIFIED NONOPIOID ANALGESIC, ANTIPYRETIC AND ANTIRHEUMATIC, INTENTIONAL SELF-HARM, SEQUELA|POISN BY UNSP NONOPI ANALGS/ANTIPYR/ANTIRHEU, SLF-HRM, SQLA
C2837947|T191|C34.00|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED MAIN BRONCHUS|MALIGNANT NEOPLASM OF UNSPECIFIED MAIN BRONCHUS
C2884800|T037|T58.8X2A|ICD10CM|TOXIC EFFECT OF CARBON MONOXIDE FROM OTHER SOURCE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CARB MONX FROM OTH SOURCE, SELF-HARM, INIT
C2884835|T037|T59.0X2S|ICD10CM|TOXIC EFFECT OF NITROGEN OXIDES, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF NITROGEN OXIDES, SELF-HARM, SEQUELA
C2838654|T037|S34.114D|ICD10CM|COMPLETE LESION OF L4 LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION OF L4 LEVEL OF LUMBAR SPINAL CORD, SUBS
C2838653|T037|S34.114A|ICD10CM|COMPLETE LESION OF L4 LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION OF L4 LEVEL OF LUMBAR SPINAL CORD, INIT
C2977856|T037|S32.509B|ICD10CM|UNSPECIFIED FRACTURE OF UNSPECIFIED PUBIS, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF UNSP PUBIS, INIT ENCNTR FOR OPEN FRACTURE
C0393819|T047|G61.81|ICD10CM|CHRONIC INFLAMMATORY DEMYELINATING POLYNEURITIS|CHRONIC INFLAMMATORY DEMYELINATING POLYNEURITIS
C0750901|T047|F00.0|DMDICD10|ALZHEIMER'S DISEASE WITH EARLY ONSET|DEMENZ BEI ALZHEIMER-KRANKHEIT, MIT FRUEHEM BEGINN (TYP 2)
C0494463|T048|F00.1|DMDICD10|ALZHEIMER'S DISEASE WITH LATE ONSET|DEMENZ BEI ALZHEIMER-KRANKHEIT, MIT SPAETEM BEGINN (TYP 1)
C0178272|T047|I28.9|DMDICD10|DISEASE OF PULMONARY VESSELS, UNSPECIFIED|KRANKHEIT DER LUNGENGEFAESSE, NICHT NAEHER BEZEICHNET
C1405840|T047||ICD10CM|OTHER DISEASES OF PULMONARY VESSELS
C0477364|T048|G30.8|DMDICD10|OTHER ALZHEIMER'S DISEASE|SONSTIGE ALZHEIMER-KRANKHEIT
C0002395|T047|G30.9|DMDICD10|ALZHEIMER'S DISEASE, UNSPECIFIED|ALZHEIMER-KRANKHEIT, NICHT NAEHER BEZEICHNET
C0155676|T046|I28.1|DMDICD10|ANEURYSM OF PULMONARY ARTERY|ANEURYSMA DER A. PULMONALIS
C0155675|T047|I28.0|DMDICD10|ARTERIOVENOUS FISTULA OF PULMONARY VESSELS|ARTERIOVENOESE FISTEL DER LUNGENGEFAESSE
C2859164|T037|S73.011A|ICD10CM|POSTERIOR SUBLUXATION OF RIGHT HIP, INITIAL ENCOUNTER|POSTERIOR SUBLUXATION OF RIGHT HIP, INITIAL ENCOUNTER
C4268130|T047|E13.3292|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|OTH DIAB WITH MILD NONP RTNOP WITHOUT MACULAR EDEMA, L EYE
C4268131|T047|E13.3293|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|OTH DIABETES WITH MILD NONP RTNOP WITHOUT MACULAR EDEMA, BI
C4268129|T047|E13.3291|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|OTH DIAB WITH MILD NONP RTNOP WITHOUT MACULAR EDEMA, R EYE
C2878586|T037|T43.612A|ICD10CM|POISONING BY CAFFEINE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY CAFFEINE, INTENTIONAL SELF-HARM, INIT ENCNTR
C4268132|T047|E13.3299|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|OTH DIAB WITH MILD NONP RTNOP WITHOUT MACULAR EDEMA, UNSP
C4268069|T047|E11.3212|ICD10CM|TYPE 2 DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|TYPE 2 DIAB WITH MILD NONP RTNOP WITH MACULAR EDEMA, L EYE
C2886087|T037|T65.4X2S|ICD10CM|TOXIC EFFECT OF CARBON DISULFIDE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CARBON DISULFIDE, SELF-HARM, SEQUELA
C4269293|T037|S02.11CA|ICD10CM|TYPE II OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE II OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, INIT
C2886104|T037|T65.5X2S|ICD10CM|TOXIC EFFECT OF NITROGLYCERIN AND OTHER NITRIC ACIDS AND ESTERS, INTENTIONAL SELF-HARM, SEQUELA|TOX EFF OF NITRO & OTH NITRIC ACIDS & ESTERS, SLF-HRM, SQLA
C4269294|T037|S02.11CB|ICD10CM|TYPE II OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE II OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, 7THB
C4267839|T191|C81.10|ICD10CM|NODULAR SCLEROSIS HODGKIN LYMPHOMA, UNSPECIFIED SITE|NODULAR SCLEROSIS HODGKIN LYMPHOMA, UNSPECIFIED SITE
C0153760|T191|C81.11|ICD10CM|NODULAR SCLEROSIS HODGKIN LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK|NODULAR SCLER HODGKIN LYMPH, NODES OF HEAD, FACE, AND NECK
C4267840|T191|C81.12|ICD10CM|NODULAR SCLEROSIS HODGKIN LYMPHOMA, INTRATHORACIC LYMPH NODES|NODULAR SCLEROSIS HODGKIN LYMPHOMA, INTRATHORAC LYMPH NODES
C4267841|T191|C81.13|ICD10CM|NODULAR SCLEROSIS HODGKIN LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES|NODULAR SCLEROSIS HODGKIN LYMPHOMA, INTRA-ABD LYMPH NODES
C0153763|T191|C81.14|ICD10CM|NODULAR SCLEROSIS HODGKIN LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB|NODULAR SCLER HODGKIN LYMPH, NODES OF AXILLA AND UPPER LIMB
C0153764|T191|C81.15|ICD10CM|NODULAR SCLEROSIS HODGKIN LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|NODLR SCLER HDGKN LYMPH, NODES OF ING REGION AND LOWER LIMB
C4267842|T191|C81.16|ICD10CM|NODULAR SCLEROSIS HODGKIN LYMPHOMA, INTRAPELVIC LYMPH NODES|NODULAR SCLEROSIS HODGKIN LYMPHOMA, INTRAPELVIC LYMPH NODES
C2018758|T191||ICD10CM|NODULAR SCLEROSIS HODGKIN LYMPHOMA, SPLEEN
C4267843|T191|C81.18|ICD10CM|NODULAR SCLEROSIS HODGKIN LYMPHOMA, LYMPH NODES OF MULTIPLE SITES|NODULAR SCLEROSIS HODGKIN LYMPHOMA, LYMPH NODES MULT SITE
C4267844|T191|C81.19|ICD10CM|NODULAR SCLEROSIS HODGKIN LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES|NODULAR SCLER HODGKIN LYMPH, EXTRNOD AND SOLID ORGAN SITES
C2886102|T037|T65.5X2A|ICD10CM|TOXIC EFFECT OF NITROGLYCERIN AND OTHER NITRIC ACIDS AND ESTERS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOX EFF OF NITRO & OTH NITRIC ACIDS & ESTERS, SLF-HRM, INIT
C4237037|T048|F12.988|ICD10CM|CANNABIS USE, UNSPECIFIED WITH OTHER CANNABIS-INDUCED DISORDER|CANNABIS INDUCED SLEEP DISORDER, WITHOUT USE DISORDER
C2853969|T191|C84.49|ICD10CM|PERIPHERAL T-CELL LYMPHOMA, NOT CLASSIFIED, EXTRANODAL AND SOLID ORGAN SITES|PRPH T-CELL LYMPH, NOT CLASS, EXTRNOD AND SOLID ORGAN SITES
C2861595|T191||ICD10CM|ACUTE PROMYELOCYTIC LEUKEMIA, IN RELAPSE
C0836971|T191||ICD10AM|ACUTE PROMYELOCYTIC LEUKEMIA, IN REMISSION
C2861594|T191||ICD10CM|ACUTE PROMYELOCYTIC LEUKEMIA, NOT HAVING ACHIEVED REMISSION
C2888818|T047|M00.062|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, LEFT KNEE|STAPHYLOCOCCAL ARTHRITIS, LEFT KNEE
C2888817|T047|M00.061|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, RIGHT KNEE|STAPHYLOCOCCAL ARTHRITIS, RIGHT KNEE
C2888819|T047|M00.069|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, UNSPECIFIED KNEE|STAPHYLOCOCCAL ARTHRITIS, UNSPECIFIED KNEE
C2874612|T048|F14.929|ICD10CM|COCAINE USE, UNSPECIFIED WITH INTOXICATION, UNSPECIFIED|COCAINE USE, UNSPECIFIED WITH INTOXICATION, UNSPECIFIED
C2873782|T047|D65|ICD10CM|DISSEMINATED INTRAVASCULAR COAGULATION [DEFIBRINATION SYNDROME]|DIFFUSE OR DISSEMINATED INTRAVASCULAR COAGULATION [DIC]
C2884366|T037|T54.1X2A|ICD10CM|TOXIC EFFECT OF OTHER CORROSIVE ORGANIC COMPOUNDS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CORROSIVE ORGANIC COMPOUNDS, SELF-HARM, INIT
C2873784|T047|D67|ICD10CM|HEREDITARY FACTOR IX DEFICIENCY|FACTOR IX DEFICIENCY (WITH FUNCTIONAL DEFECT)
C3494187|T047|D66|DMDICD10|HEREDITARY FACTOR VIII DEFICIENCY|HEREDITAERER FAKTOR-VIII-MANGEL
C2874611|T048|F14.922|ICD10CM|COCAINE USE, UNSPECIFIED WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE|COCAINE USE, UNSP W INTOXICATION WITH PERCEPTUAL DISTURBANCE
C2833585|T037|S12.600B|ICD10CM|UNSPECIFIED DISPLACED FRACTURE OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP DISP FX OF SEVENTH CERVICAL VERTEBRA, INIT FOR OPN FX
C2874609|T048|F14.920|ICD10CM|COCAINE USE, UNSPECIFIED WITH INTOXICATION, UNCOMPLICATED|COCAINE USE, UNSPECIFIED WITH INTOXICATION, UNCOMPLICATED
C2874610|T048|F14.921|ICD10CM|COCAINE USE, UNSPECIFIED WITH INTOXICATION DELIRIUM|COCAINE USE, UNSPECIFIED WITH INTOXICATION DELIRIUM
C2876895|T037|T37.4X2S|ICD10CM|POISONING BY ANTHELMINTHICS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ANTHELMINTHICS, INTENTIONAL SELF-HARM, SEQUELA
C2882805|T047|I70.408|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES, OTHER EXTREMITY|UNSP ATHSCL AUTOL VEIN BYPASS OF THE EXTRM, OTH EXTREMITY
C2882806|T047|I70.409|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES, UNSPECIFIED EXTREMITY|UNSP ATHSCL AUTOL VEIN BYPASS OF THE EXTRM, UNSP EXTREMITY
C2882803|T047|I70.402|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES, LEFT LEG|UNSP ATHSCL AUTOLOGOUS VEIN BYPASS OF THE EXTRM, LEFT LEG
C2882804|T047|I70.403|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES, BILATERAL LEGS|UNSP ATHSCL AUTOL VEIN BYPASS OF THE EXTRM, BILATERAL LEGS
C2884611|T037|T56.892S|ICD10CM|TOXIC EFFECT OF OTHER METALS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF OTHER METALS, INTENTIONAL SELF-HARM, SEQUELA
C2882802|T047|I70.401|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES, RIGHT LEG|UNSP ATHSCL AUTOLOGOUS VEIN BYPASS OF THE EXTRM, RIGHT LEG
C4268264|T048|F16.14|ICD10CM|HALLUCINOGEN ABUSE WITH HALLUCINOGEN-INDUCED MOOD DISORDER|PHENCYCLIDINE USE DISORDER, MILD, WITH PHENCYCLIDINE INDUCED DEPRESSIVE DISORDER
C4268217|T048|F12.188|ICD10CM|CANNABIS ABUSE WITH OTHER CANNABIS-INDUCED DISORDER|CANNABIS USE DISORDER, MILD, WITH CANNABIS-INDUCED SLEEP DISORDER
C2874692|T048|F16.19|ICD10CM|HALLUCINOGEN ABUSE WITH UNSPECIFIED HALLUCINOGEN-INDUCED DISORDER|HALLUCINOGEN ABUSE WITH UNSP HALLUCINOGEN-INDUCED DISORDER
C2838479|T037|S32.692A|ICD10CM|OTHER SPECIFIED FRACTURE OF LEFT ISCHIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF LEFT ISCHIUM, INIT FOR CLOS FX
C2884609|T037|T56.892A|ICD10CM|TOXIC EFFECT OF OTHER METALS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF OTH METALS, INTENTIONAL SELF-HARM, INIT
C2874481|T048|F12.180|ICD10CM|CANNABIS ABUSE WITH CANNABIS-INDUCED ANXIETY DISORDER|CANNABIS ABUSE WITH CANNABIS-INDUCED ANXIETY DISORDER
C2835797|T037|S24.131A|ICD10CM|ANTERIOR CORD SYNDROME AT T1 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|ANTERIOR CORD SYNDROME AT T1, INIT
C2890850|T037|T84.615A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL FIXATION DEVICE OF LEFT ULNA, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INT FIX OF LEFT ULNA, INIT
C0524910|T047|B18.2|DMDICD10|CHRONIC VIRAL HEPATITIS C|CHRONISCHE VIRUSHEPATITIS C
C2911652|T033|B18.1|ICD10CM|CHRONIC VIRAL HEPATITIS B WITHOUT DELTA-AGENT|CARRIER OF VIRAL HEPATITIS B
C0400918|T047|B18.0|DMDICD10|CHRONIC VIRAL HEPATITIS B WITH DELTA-AGENT|CHRONISCHE VIRUSHEPATITIS B MIT DELTA-VIRUS
C0477311|T047|D60.8|DMDICD10|OTHER ACQUIRED PURE RED CELL APLASIAS|SONSTIGE ERWORBENE ISOLIERTE APLASTISCHE ANAEMIEN
C0340961|T047|D60|DMDICD10|ACQUIRED PURE RED CELL APLASIA, UNSPECIFIED|ERWORBENE ISOLIERTE APLASTISCHE ANAEMIE [ERYTHROBLASTOPENIE] [PURE RED CELL APLASIA]
C0154043|T191|D35.4|DMDICD10|BENIGN NEOPLASM OF PINEAL GLAND|GUTARTIGE NEUBILDUNG: EPIPHYSE [GLANDULA PINEALIS] [ZIRBELDRUESE]
C0549126|T033|B18|ICD10CM|CHRONIC VIRAL HEPATITIS, UNSPECIFIED|CARRIER OF VIRAL HEPATITIS
C4267831|T033|B18.8|ICD10CM|OTHER CHRONIC VIRAL HEPATITIS|CARRIER OF OTHER VIRAL HEPATITIS
C0496901|T191|D35.2|DMDICD10|BENIGN NEOPLASM OF PITUITARY GLAND|GUTARTIGE NEUBILDUNG: HYPOPHYSE
C0451688|T047|D60.1|DMDICD10|TRANSIENT ACQUIRED PURE RED CELL APLASIA|TRANSITORISCHE ERWORBENE ISOLIERTE APLASTISCHE ANAEMIE
C4269363|T037|S02.401A|ICD10CM|MAXILLARY FRACTURE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|MAXILLARY FRACTURE, UNSPECIFIED SIDE, INIT
C4269364|T037|S02.401B|ICD10CM|MAXILLARY FRACTURE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|MAXILLARY FRACTURE, UNSPECIFIED SIDE, 7THB
C2884675|T037|T57.2X2S|ICD10CM|TOXIC EFFECT OF MANGANESE AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF MANGANESE AND ITS COMPND, SELF-HARM, SEQUELA
C2889958|T037|T82.390A|ICD10CM|OTHER MECHANICAL COMPLICATION OF AORTIC (BIFURCATION) GRAFT (REPLACEMENT), INITIAL ENCOUNTER|MECH COMPL OF AORTIC (BIFURCATION) GRAFT (REPLACEMENT), INIT
C2832411|T037|S06.386A|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF BRAINSTEM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|CONTUS/LAC/HEM BRNST W LOC >24 HR W/O RET CONSC W SURV, INIT
C4269539|T037|S02.652B|ICD10CM|FRACTURE OF ANGLE OF LEFT MANDIBLE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF ANGLE OF LEFT MANDIBLE, 7THB
C4269538|T037|S02.652A|ICD10CM|FRACTURE OF ANGLE OF LEFT MANDIBLE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF ANGLE OF LEFT MANDIBLE, INIT
C2893638|T047|M12.032|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], LEFT WRIST|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], LEFT WRIST
C2901811|T047|M86.159|ICD10CM|OTHER ACUTE OSTEOMYELITIS, UNSPECIFIED FEMUR|OTHER ACUTE OSTEOMYELITIS, UNSPECIFIED FEMUR
C2884673|T037|T57.2X2A|ICD10CM|TOXIC EFFECT OF MANGANESE AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF MANGANESE AND ITS COMPOUNDS, SELF-HARM, INIT
C2893637|T047|M12.031|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], RIGHT WRIST|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], RIGHT WRIST
C2901809|T047|M86.151|ICD10CM|OTHER ACUTE OSTEOMYELITIS, RIGHT FEMUR|OTHER ACUTE OSTEOMYELITIS, RIGHT FEMUR
C2832413|T037|S06.386S|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF BRAINSTEM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|CONTUS/LAC/HEM BRNST W LOC >24 HR W/O RET CONSC W SURV, SQLA
C2901810|T047|M86.152|ICD10CM|OTHER ACUTE OSTEOMYELITIS, LEFT FEMUR|OTHER ACUTE OSTEOMYELITIS, LEFT FEMUR
C2889275|T047|M05.532|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT WRIST|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF LEFT WRIST
C0268583|T047|E71.120|ICD10CM|METHYLMALONIC ACIDEMIA|METHYLMALONIC ACIDEMIA
C2889274|T047|M05.531|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT WRIST|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT WRIST
C2874238|T047|E71.128|ICD10CM|OTHER DISORDERS OF PROPIONATE METABOLISM|OTHER DISORDERS OF PROPIONATE METABOLISM
C2889276|T047|M05.539|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP WRIST
C2835306|T037|S22.041B|ICD10CM|STABLE BURST FRACTURE OF FOURTH THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|STABLE BURST FX FOURTH THOR VERTEBRA, INIT FOR OPN FX
C2835305|T037|S22.041A|ICD10CM|STABLE BURST FRACTURE OF FOURTH THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|STABLE BURST FRACTURE OF FOURTH THORACIC VERTEBRA, INIT
C3264223|T047|H40.1332|ICD10CM|PIGMENTARY GLAUCOMA, BILATERAL, MODERATE STAGE|PIGMENTARY GLAUCOMA, BILATERAL, MODERATE STAGE
C3264224|T047|H40.1333|ICD10CM|PIGMENTARY GLAUCOMA, BILATERAL, SEVERE STAGE|PIGMENTARY GLAUCOMA, BILATERAL, SEVERE STAGE
C3264221|T047|H40.1330|ICD10CM|PIGMENTARY GLAUCOMA, BILATERAL, STAGE UNSPECIFIED|PIGMENTARY GLAUCOMA, BILATERAL, STAGE UNSPECIFIED
C3264222|T047|H40.1331|ICD10CM|PIGMENTARY GLAUCOMA, BILATERAL, MILD STAGE|PIGMENTARY GLAUCOMA, BILATERAL, MILD STAGE
C4290157|T047|I70.35|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF OTHER EXTREMITY WITH ULCERATION|ANY CONDITION CLASSIFIABLE TO I70.318 AND I70.328
C3264225|T047|H40.1334|ICD10CM|PIGMENTARY GLAUCOMA, BILATERAL, INDETERMINATE STAGE|PIGMENTARY GLAUCOMA, BILATERAL, INDETERMINATE STAGE
C2889326|T047|M05.70|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED SITE WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRITIS W RHEU FACTOR OF UNSP SITE W/O ORG/SYS INVOLV
C2889355|T047|M05.79|ICD10CM|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF MULTIPLE SITES WITHOUT ORGAN OR SYSTEMS INVOLVEMENT|RHEU ARTHRITIS W RHEU FACTOR MULT SITE W/O ORG/SYS INVOLV
C2874769|T048|F18.280|ICD10CM|INHALANT DEPENDENCE WITH INHALANT-INDUCED ANXIETY DISORDER|INHALANT DEPENDENCE WITH INHALANT-INDUCED ANXIETY DISORDER
C4268095|T047|E11.3519|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|TYPE 2 DIAB WITH PROLIF DIAB RTNOP WITH MACULAR EDEMA, UNSP
C4268094|T047|E11.3513|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|TYPE 2 DIAB WITH PROLIF DIAB RTNOP WITH MACULAR EDEMA, BI
C4268093|T047|E11.3512|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|TYPE 2 DIAB WITH PROLIF DIAB RTNOP WITH MACULAR EDEMA, L EYE
C4268092|T047|E11.3511|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|TYPE 2 DIAB WITH PROLIF DIAB RTNOP WITH MACULAR EDEMA, R EYE
C4268414|T047|H40.1194|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, UNSPECIFIED EYE, INDETERMINATE STAGE|PRIMARY OPEN-ANGLE GLAUCOMA, UNSP, INDETERMINATE STAGE
C2874373|T048|F10.121|ICD10CM|ALCOHOL ABUSE WITH INTOXICATION DELIRIUM|ALCOHOL ABUSE WITH INTOXICATION DELIRIUM
C4268412|T047|H40.1192|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, UNSPECIFIED EYE, MODERATE STAGE|PRIMARY OPEN-ANGLE GLAUCOMA, UNSPECIFIED EYE, MODERATE STAGE
C4268413|T047|H40.1193|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, UNSPECIFIED EYE, SEVERE STAGE|PRIMARY OPEN-ANGLE GLAUCOMA, UNSPECIFIED EYE, SEVERE STAGE
C4268410|T047|H40.1190|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, UNSPECIFIED EYE, STAGE UNSPECIFIED|PRIMARY OPEN-ANGLE GLAUCOMA, UNSP, STAGE UNSPECIFIED
C4268411|T047|H40.1191|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, UNSPECIFIED EYE, MILD STAGE|PRIMARY OPEN-ANGLE GLAUCOMA, UNSPECIFIED EYE, MILD STAGE
C2858544|T037|S72.431C|ICD10CM|DISPLACED FRACTURE OF MEDIAL CONDYLE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF MED CONDYLE OF R FEMR, 7THC
C2858543|T037|S72.431B|ICD10CM|DISPLACED FRACTURE OF MEDIAL CONDYLE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF MED CONDYLE OF R FEMUR, INIT FOR OPN FX TYPE I/2
C2858542|T037|S72.431A|ICD10CM|DISPLACED FRACTURE OF MEDIAL CONDYLE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF MEDIAL CONDYLE OF RIGHT FEMUR, INIT FOR CLOS FX
C2874371|T048|F10.129|ICD10CM|ALCOHOL ABUSE WITH INTOXICATION, UNSPECIFIED|ALCOHOL ABUSE WITH INTOXICATION, UNSPECIFIED
C2834033|T037|S14.151D|ICD10CM|OTHER INCOMPLETE LESION AT C1 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|OTH INCOMPLETE LESION AT C1, SUBS
C2834034|T037|S14.151S|ICD10CM|OTHER INCOMPLETE LESION AT C1 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|OTH INCOMPLETE LESION AT C1, SEQUELA
C2905688|T037|X73.8XXD|ICD10CM|INTENTIONAL SELF-HARM BY OTHER LARGER FIREARM DISCHARGE, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY OTH LARGER FIREARM DISCHARGE, SUBS
C2843286|T037|S48.022A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEFT SHOULDER JOINT, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION AT LEFT SHOULDER JOINT, INIT
C2856812|T037|S72.042C|ICD10CM|DISPLACED FRACTURE OF BASE OF NECK OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF BASE OF NK OF L FEMR, INIT FOR OPN FX TYPE 3A/B/C
C2843288|T037|S48.022S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEFT SHOULDER JOINT, SEQUELA|PARTIAL TRAUMATIC AMPUTATION AT LEFT SHOULDER JOINT, SEQUELA
C2859177|T037|S73.015A|ICD10CM|POSTERIOR DISLOCATION OF LEFT HIP, INITIAL ENCOUNTER|POSTERIOR DISLOCATION OF LEFT HIP, INITIAL ENCOUNTER
C2834018|T037|S14.147D|ICD10CM|BROWN-SEQUARD SYNDROME AT C7 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|BROWN-SEQUARD SYNDROME AT C7, SUBS
C0155764|T047|I77.9|DMDICD10|DISORDER OF ARTERIES AND ARTERIOLES, UNSPECIFIED|KRANKHEIT DER ARTERIEN UND ARTERIOLEN, NICHT NAEHER BEZEICHNET
C0155762|T047|I77.5|DMDICD10|NECROSIS OF ARTERY|ARTERIENNEKROSE
C1861783|T047|I77.4|DMDICD10|CELIAC ARTERY COMPRESSION SYNDROME|ARTERIA-COELIACA-KOMPRESSIONS-SYNDROM
C0014100|T047||ICD10CM|ARTERITIS, UNSPECIFIED
C1388472|T190||ICD10CM|STRICTURE OF ARTERY
C1541850|T020|I77.0|DMDICD10|ARTERIOVENOUS FISTULA, ACQUIRED|ARTERIOVENOESE FISTEL, ERWORBEN
C1998294|T047||ICD10CM|ARTERIAL FIBROMUSCULAR DYSPLASIA
C0265000|T047|I77.2|ICD10CM|RUPTURE OF ARTERY|ULCER OF ARTERY
C2842132|T191|C50.822|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF LEFT MALE BREAST|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF LEFT MALE BREAST
C0494675|T047|J69.1|DMDICD10|PNEUMONITIS DUE TO INHALATION OF OILS AND ESSENCES|PNEUMONIE DURCH OELE UND EXTRAKTE
C2887481|T047|J69.0|ICD10CM|PNEUMONITIS DUE TO INHALATION OF FOOD AND VOMIT|PNEUMONITIS DUE TO INHALATION OF FOOD AND VOMIT
C2890509|T037|T84.051A|ICD10CM|PERIPROSTHETIC OSTEOLYSIS OF INTERNAL PROSTHETIC LEFT HIP JOINT, INITIAL ENCOUNTER|PERIPROSTH OSTEOLYSIS OF INTERNAL PROSTHETIC L HIP JT, INIT
C2887483|T037|J69.8|ICD10CM|PNEUMONITIS DUE TO INHALATION OF OTHER SOLIDS AND LIQUIDS|PNEUMONITIS DUE TO ASPIRATION OF DETERGENT
C2902105|T046|M87.350|ICD10CM|OTHER SECONDARY OSTEONECROSIS, PELVIS|OTHER SECONDARY OSTEONECROSIS, PELVIS
C2902106|T046|M87.351|ICD10CM|OTHER SECONDARY OSTEONECROSIS, RIGHT FEMUR|OTHER SECONDARY OSTEONECROSIS, RIGHT FEMUR
C2902107|T046|M87.352|ICD10CM|OTHER SECONDARY OSTEONECROSIS, LEFT FEMUR|OTHER SECONDARY OSTEONECROSIS, LEFT FEMUR
C2902108|T046|M87.353|ICD10CM|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED FEMUR|OTHER SECONDARY OSTEONECROSIS, UNSPECIFIED FEMUR
C4268053|T047|E10.3549|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, UNSPECIFIED EYE|TYPE 1 DIAB WITH PROLIF DIAB RTNOP WITH COMB DETACH, UNSP
C2857856|T037|S72.333A|ICD10CM|DISPLACED OBLIQUE FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED OBLIQUE FRACTURE OF SHAFT OF UNSP FEMUR, INIT
C2857857|T037|S72.333B|ICD10CM|DISPLACED OBLIQUE FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL OBLIQUE FX SHAFT OF UNSP FEMR, 7THB
C2857858|T037|S72.333C|ICD10CM|DISPLACED OBLIQUE FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL OBLIQUE FX SHAFT OF UNSP FEMR, 7THC
C2890720|T037|T84.226A|ICD10CM|DISPLACEMENT OF INTERNAL FIXATION DEVICE OF VERTEBRAE, INITIAL ENCOUNTER|DISPLACEMENT OF INTERNAL FIXATION DEVICE OF VERTEBRAE, INIT
C2901574|T046|M84.675A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, LEFT FOOT, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, LEFT FOOT, INIT FOR FX
C2896684|T046|M80.821A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, RIGHT HUMERUS, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, R HUMERUS, INIT
C2883026|T047|I70.798|ICD10CM|OTHER ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, OTHER EXTREMITY|OTH ATHSCL TYPE OF BYPASS OF THE EXTREMITIES, OTH EXTREMITY
C2883027|T047|I70.799|ICD10CM|OTHER ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, UNSPECIFIED EXTREMITY|OTH ATHSCL TYPE OF BYPASS OF THE EXTREMITIES, UNSP EXTREMITY
C2883024|T047|I70.792|ICD10CM|OTHER ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, LEFT LEG|OTH ATHSCL TYPE OF BYPASS OF THE EXTREMITIES, LEFT LEG
C2883025|T047|I70.793|ICD10CM|OTHER ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, BILATERAL LEGS|OTH ATHSCL TYPE OF BYPASS OF THE EXTREMITIES, BILATERAL LEGS
C2883023|T047|I70.791|ICD10CM|OTHER ATHEROSCLEROSIS OF OTHER TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, RIGHT LEG|OTH ATHSCL TYPE OF BYPASS OF THE EXTREMITIES, RIGHT LEG
C2888904|T047|M00.831|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, RIGHT WRIST|ARTHRITIS DUE TO OTHER BACTERIA, RIGHT WRIST
C2888905|T047|M00.832|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, LEFT WRIST|ARTHRITIS DUE TO OTHER BACTERIA, LEFT WRIST
C3161078|T048|F03.90|ICD10CM|UNSPECIFIED DEMENTIA WITHOUT BEHAVIORAL DISTURBANCE|UNSPECIFIED DEMENTIA WITHOUT BEHAVIORAL DISTURBANCE
C2890243|T037|T83.110A|ICD10CM|BREAKDOWN (MECHANICAL) OF URINARY ELECTRONIC STIMULATOR DEVICE, INITIAL ENCOUNTER|BREAKDOWN OF URINARY ELECTRONIC STIMULATOR DEVICE, INIT
C2888906|T047|M00.839|ICD10CM|ARTHRITIS DUE TO OTHER BACTERIA, UNSPECIFIED WRIST|ARTHRITIS DUE TO OTHER BACTERIA, UNSPECIFIED WRIST
C2939420|T191||ICD10CM|SECONDARY MALIGNANT NEOPLASM OF UNSPECIFIED SITE
C0153349|T191|C02.9|DMDICD10|MALIGNANT NEOPLASM OF TONGUE, UNSPECIFIED|BOESARTIGE NEUBILDUNG: ZUNGE, NICHT NAEHER BEZEICHNET
C2833835|T191|C02.8|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF TONGUE|MALIGNANT NEOPLASM OF TWO OR MORE CONTIGUOUS SITES OF TONGUE
C0153356|T191|C02.4|DMDICD10|MALIGNANT NEOPLASM OF LINGUAL TONSIL|BOESARTIGE NEUBILDUNG: ZUNGENTONSILLE
C2833834|T191|C02.3|ICD10CM|MALIGNANT NEOPLASM OF ANTERIOR TWO-THIRDS OF TONGUE, PART UNSPECIFIED|MALIGNANT NEOPLASM OF MIDDLE THIRD OF TONGUE NOS
C0684333|T191|C02.2|DMDICD10|MALIGNANT NEOPLASM OF VENTRAL SURFACE OF TONGUE|BOESARTIGE NEUBILDUNG: ZUNGENUNTERFLAECHE
C0496755|T191|C02.1|DMDICD10|MALIGNANT NEOPLASM OF BORDER OF TONGUE|BOESARTIGE NEUBILDUNG: ZUNGENRAND
C2521535|T060|C020|ICD10PCS|MALIGNANT NEOPLASM OF DORSAL SURFACE OF TONGUE|NUCLEAR MEDICINE @ CENTRAL NERVOUS SYSTEM @ TOMOGRAPHIC (TOMO) NUCLEAR MEDICINE IMAGING @ BRAIN
C2838344|T037|S32.486B|ICD10CM|NONDISPLACED DOME FRACTURE OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP DOME FRACTURE OF UNSP ACETABULUM, INIT FOR OPN FX
C2889923|T037|T82.322A|ICD10CM|DISPLACEMENT OF FEMORAL ARTERIAL GRAFT (BYPASS), INITIAL ENCOUNTER|DISPLACEMENT OF FEMORAL ARTERIAL GRAFT (BYPASS), INIT ENCNTR
C4269489|T037|S02.631A|ICD10CM|FRACTURE OF CORONOID PROCESS OF RIGHT MANDIBLE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF CORONOID PROCESS OF RIGHT MANDIBLE, INIT
C4269490|T037|S02.631B|ICD10CM|FRACTURE OF CORONOID PROCESS OF RIGHT MANDIBLE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF CORONOID PROCESS OF RIGHT MANDIBLE, 7THB
C2876796|T037|T37.0X2S|ICD10CM|POISONING BY SULFONAMIDES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY SULFONAMIDES, INTENTIONAL SELF-HARM, SEQUELA
C0750952|T191|C24.9|DMDICD10|MALIGNANT NEOPLASM OF BILIARY TRACT, UNSPECIFIED|BOESARTIGE NEUBILDUNG: GALLENWEGE, NICHT NAEHER BEZEICHNET
C2837939|T191|C24.8|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF BILIARY TRACT|PRIMARY MALIGNANT NEOPLASM OF TWO OR MORE CONTIGUOUS SITES OF BILIARY TRACT
C0153454|T191|C24.1|DMDICD10|MALIGNANT NEOPLASM OF AMPULLA OF VATER|BOESARTIGE NEUBILDUNG: AMPULLA HEPATOPANCREATICA [AMPULLA VATERI]
C3665467|T191|C24.0|ICD10CM|MALIGNANT NEOPLASM OF EXTRAHEPATIC BILE DUCT|MALIGNANT NEOPLASM OF COMMON BILE DUCT
C4270280|T046|T83.24XA|ICD10CM|EROSION OF GRAFT OF URINARY ORGAN, INITIAL ENCOUNTER|EROSION OF GRAFT OF URINARY ORGAN, INITIAL ENCOUNTER
C1399675|T047||ICD10CM|HEMOPHAGOCYTIC LYMPHOHISTIOCYTOSIS
C2832056|T037|S06.300S|ICD10CM|UNSPECIFIED FOCAL TRAUMATIC BRAIN INJURY WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|UNSP FOCAL TBI W/O LOSS OF CONSCIOUSNESS, SEQUELA
C2874815|T048|F19.22|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH INTOXICATION, UNSPECIFIED|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH INTOXICATION
C2837736|T037|S32.131A|ICD10CM|MINIMALLY DISPLACED ZONE III FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|MINIMALLY DISPLACED ZONE III FRACTURE OF SACRUM, INIT
C2832054|T037|S06.300A|ICD10CM|UNSPECIFIED FOCAL TRAUMATIC BRAIN INJURY WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|UNSP FOCAL TBI W/O LOSS OF CONSCIOUSNESS, INIT
C2745961|T191|C78.39|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF OTHER RESPIRATORY ORGANS|SECONDARY MALIGNANT NEOPLASM OF OTHER RESPIRATORY ORGANS
C2888576|T047|L89.624|ICD10CM|PRESSURE ULCER OF LEFT HEEL, STAGE 4|PRESSURE ULCER OF LEFT HEEL, STAGE 4
C2845960|T191|C78.30|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF UNSPECIFIED RESPIRATORY ORGAN|SECONDARY MALIGNANT NEOPLASM OF UNSP RESPIRATORY ORGAN
C2885966|T037|T64.82XA|ICD10CM|TOXIC EFFECT OF OTHER MYCOTOXIN FOOD CONTAMINANTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF MYCOTOXIN FOOD CONTAMINANTS, SELF-HARM, INIT
C2856637|T037|S72.024A|ICD10CM|NONDISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF EPIPHY (SEPARATION) (UPPER) OF R FEMUR, INIT
C2885711|T037|T63.482A|ICD10CM|TOXIC EFFECT OF VENOM OF OTHER ARTHROPOD, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF ARTHROPOD, SELF-HARM, INIT
C2882276|T047|I50.43|ICD10CM|ACUTE ON CHRONIC COMBINED SYSTOLIC (CONGESTIVE) AND DIASTOLIC (CONGESTIVE) HEART FAILURE|ACUTE ON CHRONIC COMBINED SYSTOLIC (CONGESTIVE) AND DIASTOLIC (CONGESTIVE) HEART FAILURE
C2882275|T047|I50.42|ICD10CM|CHRONIC COMBINED SYSTOLIC (CONGESTIVE) AND DIASTOLIC (CONGESTIVE) HEART FAILURE|CHRONIC COMBINED SYSTOLIC (CONGESTIVE) AND DIASTOLIC (CONGESTIVE) HEART FAILURE
C2882274|T047|I50.41|ICD10CM|ACUTE COMBINED SYSTOLIC (CONGESTIVE) AND DIASTOLIC (CONGESTIVE) HEART FAILURE|ACUTE COMBINED SYSTOLIC (CONGESTIVE) AND DIASTOLIC (CONGESTIVE) HEART FAILURE
C2882273|T047|I50.40|ICD10CM|UNSPECIFIED COMBINED SYSTOLIC (CONGESTIVE) AND DIASTOLIC (CONGESTIVE) HEART FAILURE|UNSP COMBINED SYSTOLIC AND DIASTOLIC (CONGESTIVE) HRT FAIL
C2885968|T037|T64.82XS|ICD10CM|TOXIC EFFECT OF OTHER MYCOTOXIN FOOD CONTAMINANTS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF MYCOTOXIN FOOD CONTAMNT, SELF-HARM, SEQUELA
C2856639|T037|S72.024C|ICD10CM|NONDISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF EPIPHY (SEPARATION) (UPPER) OF R FEMR, 7THC
C2853889|T191|C83.05|ICD10CM|SMALL CELL B-CELL LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|SMALL CELL B-CELL LYMPH, NODES OF ING REGION AND LOWER LIMB
C2853888|T191|C83.04|ICD10CM|SMALL CELL B-CELL LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB|SMALL CELL B-CELL LYMPHOMA, NODES OF AXILLA AND UPPER LIMB
C2873953|T047|E09.10|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH KETOACIDOSIS WITHOUT COMA|DRUG/CHEM DIABETES MELLITUS W KETOACIDOSIS W/O COMA
C2873954|T047|E09.11|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH KETOACIDOSIS WITH COMA|DRUG/CHEM DIABETES MELLITUS W KETOACIDOSIS W COMA
C2853885|T191|C83.01|ICD10CM|SMALL CELL B-CELL LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK|SMALL CELL B-CELL LYMPHOMA, NODES OF HEAD, FACE, AND NECK
C2853884|T191|C83.00|ICD10CM|SMALL CELL B-CELL LYMPHOMA, UNSPECIFIED SITE|SMALL CELL B-CELL LYMPHOMA, UNSPECIFIED SITE
C2853887|T191|C83.03|ICD10CM|SMALL CELL B-CELL LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES|SMALL CELL B-CELL LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES
C2853886|T191|C83.02|ICD10CM|SMALL CELL B-CELL LYMPHOMA, INTRATHORACIC LYMPH NODES|SMALL CELL B-CELL LYMPHOMA, INTRATHORACIC LYMPH NODES
C2883964|T037|T50.Z92S|ICD10CM|POISONING BY OTHER VACCINES AND BIOLOGICAL SUBSTANCES, INTENTIONAL SELF-HARM, SEQUELA|POISN BY OTH VACCINES AND BIOLG SUBSTNC, SELF-HARM, SEQUELA
C0036939|T048|F24|DMDICD10|SHARED PSYCHOTIC DISORDER|INDUZIERTE WAHNHAFTE STOERUNG
C2853893|T191|C83.09|ICD10CM|SMALL CELL B-CELL LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES|SMALL CELL B-CELL LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES
C2853892|T191|C83.08|ICD10CM|SMALL CELL B-CELL LYMPHOMA, LYMPH NODES OF MULTIPLE SITES|SMALL CELL B-CELL LYMPHOMA, LYMPH NODES OF MULTIPLE SITES
C2902901|T047|N05.6|ICD10CM|UNSPECIFIED NEPHRITIC SYNDROME WITH DENSE DEPOSIT DISEASE|UNSPECIFIED NEPHRITIC SYNDROME WITH MEMBRANOPROLIFERATIVE GLOMERULONEPHRITIS, TYPE 2
C2882658|T046|I69.931|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING RIGHT DOMINANT SIDE|MONOPLG UPR LMB FOL UNSP CEREBVASC DIS AFF RIGHT DOM SIDE
C2883962|T037|T50.Z92A|ICD10CM|POISONING BY OTHER VACCINES AND BIOLOGICAL SUBSTANCES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH VACCINES AND BIOLG SUBSTNC, SELF-HARM, INIT
C2902899|T047|N05.1|ICD10CM|UNSPECIFIED NEPHRITIC SYNDROME WITH FOCAL AND SEGMENTAL GLOMERULAR LESIONS|UNSPECIFIED NEPHRITIC SYNDROME WITH FOCAL GLOMERULONEPHRITIS
C2882659|T046|I69.932|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING LEFT DOMINANT SIDE|MONOPLG UPR LMB FOL UNSP CEREBVASC DISEASE AFF LEFT DOM SIDE
C2901372|T046|M84.611A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, RIGHT SHOULDER, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, RIGHT SHOULDER, INIT
C2880090|T047|A01.05|ICD10CM|TYPHOID OSTEOMYELITIS|TYPHOID OSTEOMYELITIS
C2882661|T046|I69.934|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING LEFT NON-DOMINANT SIDE|MONOPLG UPR LMB FOL UNSP CEREBVASC DIS AFF LEFT NONDOM SIDE
C0339956|T047|A01.03|ICD10CM|TYPHOID PNEUMONIA|TYPHOID PNEUMONIA
C2901875|T047|M86.432|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, LEFT RADIUS AND ULNA|CHRONIC OSTEOMYELITIS W DRAINING SINUS, LEFT RADIUS AND ULNA
C2901874|T047|M86.431|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, RIGHT RADIUS AND ULNA|CHRONIC OSTEOMYELIT W DRAINING SINUS, RIGHT RADIUS AND ULNA
C2901876|T047|M86.439|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, UNSPECIFIED RADIUS AND ULNA|CHRONIC OSTEOMYELITIS W DRAINING SINUS, UNSP RADIUS AND ULNA
C2833948|T037|S14.128D|ICD10CM|CENTRAL CORD SYNDROME AT C8 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|CENTRAL CORD SYNDROME AT C8, SUBS
C2838294|T037|S32.475B|ICD10CM|NONDISPLACED FRACTURE OF MEDIAL WALL OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP FX OF MEDIAL WALL OF LEFT ACETAB, INIT FOR OPN FX
C2838293|T037|S32.475A|ICD10CM|NONDISPLACED FRACTURE OF MEDIAL WALL OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF MEDIAL WALL OF LEFT ACETABULUM, INIT
C0477376|T047|G46.7|DMDICD10|OTHER LACUNAR SYNDROMES|SONSTIGE LAKUNAERE SYNDROME
C2902904|T047|N05.8|ICD10CM|UNSPECIFIED NEPHRITIC SYNDROME WITH OTHER MORPHOLOGIC CHANGES|UNSP NEPHRITIC SYNDROME WITH OTHER MORPHOLOGIC CHANGES
C2874605|T048|F14.29|ICD10CM|COCAINE DEPENDENCE WITH UNSPECIFIED COCAINE-INDUCED DISORDER|COCAINE DEPENDENCE WITH UNSPECIFIED COCAINE-INDUCED DISORDER
C0339904|T047||ICD10CM|SYSTEMIC SCLEROSIS WITH LUNG INVOLVEMENT
C2895197|T047|M34.83|ICD10CM|SYSTEMIC SCLEROSIS WITH POLYNEUROPATHY|SYSTEMIC SCLEROSIS WITH POLYNEUROPATHY
C2895196|T047|M34.82|ICD10CM|SYSTEMIC SCLEROSIS WITH MYOPATHY|SYSTEMIC SCLEROSIS WITH MYOPATHY
C2874595|T048|F14.23|ICD10CM|COCAINE DEPENDENCE WITH WITHDRAWAL|COCAINE DEPENDENCE WITH WITHDRAWAL
C4237066|T048|F14.20|ICD10CM|COCAINE DEPENDENCE, UNCOMPLICATED|COCAINE USE DISORDER, SEVERE
C4509061|T048|F14.21|ICD10CM|COCAINE DEPENDENCE, IN REMISSION|COCAINE USE DISORDER, SEVERE, IN SUSTAINED REMISSION
C2895198|T047|M34.89|ICD10CM|OTHER SYSTEMIC SCLEROSIS|OTHER SYSTEMIC SCLEROSIS
C4268238|T048|F14.24|ICD10CM|COCAINE DEPENDENCE WITH COCAINE-INDUCED MOOD DISORDER|COCAINE USE DISORDER, SEVERE, WITH COCAINE-INDUCED DEPRESSIVE DISORDER
C2855964|T037|S68.422A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT HAND AT WRIST LEVEL, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP OF LEFT HAND AT WRIST LEVEL, INIT
C2859244|T037|S73.043A|ICD10CM|CENTRAL SUBLUXATION OF UNSPECIFIED HIP, INITIAL ENCOUNTER|CENTRAL SUBLUXATION OF UNSPECIFIED HIP, INITIAL ENCOUNTER
C2888858|T047|M00.19|ICD10CM|PNEUMOCOCCAL POLYARTHRITIS|PNEUMOCOCCAL POLYARTHRITIS
C2888857|T047||ICD10CM|PNEUMOCOCCAL ARTHRITIS, VERTEBRAE
C2888827|T047|M00.10|ICD10CM|PNEUMOCOCCAL ARTHRITIS, UNSPECIFIED JOINT|PNEUMOCOCCAL ARTHRITIS, UNSPECIFIED JOINT
C3264210|T047|H40.1294|ICD10CM|LOW-TENSION GLAUCOMA, UNSPECIFIED EYE, INDETERMINATE STAGE|LOW-TENSION GLAUCOMA, UNSPECIFIED EYE, INDETERMINATE STAGE
C3264207|T047|H40.1291|ICD10CM|LOW-TENSION GLAUCOMA, UNSPECIFIED EYE, MILD STAGE|LOW-TENSION GLAUCOMA, UNSPECIFIED EYE, MILD STAGE
C3264206|T047|H40.1290|ICD10CM|LOW-TENSION GLAUCOMA, UNSPECIFIED EYE, STAGE UNSPECIFIED|LOW-TENSION GLAUCOMA, UNSPECIFIED EYE, STAGE UNSPECIFIED
C3264209|T047|H40.1293|ICD10CM|LOW-TENSION GLAUCOMA, UNSPECIFIED EYE, SEVERE STAGE|LOW-TENSION GLAUCOMA, UNSPECIFIED EYE, SEVERE STAGE
C3264208|T047|H40.1292|ICD10CM|LOW-TENSION GLAUCOMA, UNSPECIFIED EYE, MODERATE STAGE|LOW-TENSION GLAUCOMA, UNSPECIFIED EYE, MODERATE STAGE
C2889563|T047|M08.25|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, UNSPECIFIED HIP|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, HIP
C2889564|T047|M08.251|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, RIGHT HIP|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, RIGHT HIP
C2889565|T047|M08.252|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, LEFT HIP|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, LEFT HIP
C2833152|T037|S12.01XA|ICD10CM|STABLE BURST FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|STABLE BURST FRACTURE OF FIRST CERVICAL VERTEBRA, INIT
C2833153|T037|S12.01XB|ICD10CM|STABLE BURST FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|STABLE BURST FX FIRST CERVCAL VERTEBRA, INIT FOR OPN FX
C2888872|T047|M00.239|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, UNSPECIFIED WRIST|OTHER STREPTOCOCCAL ARTHRITIS, UNSPECIFIED WRIST
C2888871|T047|M00.232|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, LEFT WRIST|OTHER STREPTOCOCCAL ARTHRITIS, LEFT WRIST
C0348818|T047|J44.0|DMDICD10|CHRONIC OBSTRUCTIVE PULMONARY DISEASE WITH ACUTE LOWER RESPIRATORY INFECTION|CHRONISCHE OBSTRUKTIVE LUNGENKRANKHEIT MIT AKUTER INFEKTION DER UNTEREN ATEMWEGE
C2888870|T047|M00.231|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, RIGHT WRIST|OTHER STREPTOCOCCAL ARTHRITIS, RIGHT WRIST
C0546982|T047||ICD10CM|MECONIUM ILEUS IN CYSTIC FIBROSIS
C2874308|T047|E84.19|ICD10CM|CYSTIC FIBROSIS WITH OTHER INTESTINAL MANIFESTATIONS|CYSTIC FIBROSIS WITH OTHER INTESTINAL MANIFESTATIONS
C4270355|T046|T83.61XA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO IMPLANTED PENILE PROSTHESIS, INITIAL ENCOUNTER|I/I REACT D/T IMPLANTED PENILE PROSTHESIS, INITIAL ENCOUNTER
C2921069|T047||ICD10CM|THORACIC AORTIC ECTASIA
C2921070|T047|I77.811|ICD10CM|ABDOMINAL AORTIC ECTASIA|ABDOMINAL AORTIC ECTASIA
C2921071|T047||ICD10CM|THORACOABDOMINAL AORTIC ECTASIA
C2889532|T047|M08.031|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, RIGHT WRIST|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, RIGHT WRIST
C2889533|T047|M08.032|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, LEFT WRIST|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, LEFT WRIST
C2921068|T047|I77.819|ICD10CM|AORTIC ECTASIA, UNSPECIFIED SITE|AORTIC ECTASIA, UNSPECIFIED SITE
C2889534|T047|M08.03|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED WRIST|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, WRIST
C2876146|T037|T31.54|ICD10CM|BURNS INVOLVING 50-59% OF BODY SURFACE WITH 40-49% THIRD DEGREE BURNS|BURNS OF 50-59% OF BODY SURFACE W 40-49% THIRD DEGREE BURNS
C2876147|T037|T31.55|ICD10CM|BURNS INVOLVING 50-59% OF BODY SURFACE WITH 50-59% THIRD DEGREE BURNS|BURNS OF 50-59% OF BODY SURFACE W 50-59% THIRD DEGREE BURNS
C2876144|T037|T31.52|ICD10CM|BURNS INVOLVING 50-59% OF BODY SURFACE WITH 20-29% THIRD DEGREE BURNS|BURNS OF 50-59% OF BODY SURFACE W 20-29% THIRD DEGREE BURNS
C2876145|T037|T31.53|ICD10CM|BURNS INVOLVING 50-59% OF BODY SURFACE WITH 30-39% THIRD DEGREE BURNS|BURNS OF 50-59% OF BODY SURFACE W 30-39% THIRD DEGREE BURNS
C2876143|T037|T31.51|ICD10CM|BURNS INVOLVING 50-59% OF BODY SURFACE WITH 10-19% THIRD DEGREE BURNS|BURNS OF 50-59% OF BODY SURFACE W 10-19% THIRD DEGREE BURNS
C2832629|T037|S06.829S|ICD10CM|INJURY OF LEFT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|INJ L INT CAROTID, INTCR W LOC OF UNSP DURATION, SEQUELA
C2832627|T037|S06.829A|ICD10CM|INJURY OF LEFT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|INJURY OF L INT CAROTID, INTCR W LOC OF UNSP DURATION, INIT
C2888940|T047|M01.X39|ICD10CM|DIRECT INFECTION OF UNSPECIFIED WRIST IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIR INFCT OF UNSP WRIST IN INFEC/PARASTC DIS CLASSD ELSWHR
C2888939|T047|M01.X32|ICD10CM|DIRECT INFECTION OF LEFT WRIST IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIRECT INFCT OF L WRIST IN INFEC/PARASTC DIS CLASSD ELSWHR
C2888938|T047|M01.X31|ICD10CM|DIRECT INFECTION OF RIGHT WRIST IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIRECT INFCT OF R WRIST IN INFEC/PARASTC DIS CLASSD ELSWHR
C2890646|T037|T84.127A|ICD10CM|DISPLACEMENT OF INTERNAL FIXATION DEVICE OF BONE OF LEFT LOWER LEG, INITIAL ENCOUNTER|DISPLACEMENT OF INT FIX OF BONE OF LEFT LOWER LEG, INIT
C0840049|T046|M87.89|ICD10CM|OTHER OSTEONECROSIS, MULTIPLE SITES|OTHER OSTEONECROSIS, MULTIPLE SITES
C2902020|T046|M87.166|ICD10CM|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED FIBULA|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED FIBULA
C2902019|T046|M87.165|ICD10CM|OSTEONECROSIS DUE TO DRUGS, LEFT FIBULA|OSTEONECROSIS DUE TO DRUGS, LEFT FIBULA
C2902018|T046|M87.164|ICD10CM|OSTEONECROSIS DUE TO DRUGS, RIGHT FIBULA|OSTEONECROSIS DUE TO DRUGS, RIGHT FIBULA
C2902017|T046|M87.163|ICD10CM|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED TIBIA|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED TIBIA
C2902016|T046|M87.162|ICD10CM|OSTEONECROSIS DUE TO DRUGS, LEFT TIBIA|OSTEONECROSIS DUE TO DRUGS, LEFT TIBIA
C2902015|T046|M87.161|ICD10CM|OSTEONECROSIS DUE TO DRUGS, RIGHT TIBIA|OSTEONECROSIS DUE TO DRUGS, RIGHT TIBIA
C2887361|T047|I97.811|ICD10CM|INTRAOPERATIVE CEREBROVASCULAR INFARCTION DURING OTHER SURGERY|INTRAOPERATIVE CEREBROVASCULAR INFARCTION DURING OTH SURGERY
C2845938|T191|C72.50|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED CRANIAL NERVE|MALIGNANT NEOPLASM OF UNSPECIFIED CRANIAL NERVE
C4270615|T046|T85.820A|ICD10CM|FIBROSIS DUE TO NERVOUS SYSTEM PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|FIBROSIS DUE TO NERVOUS SYSTEM PROSTH DEV/GRFT, INIT
C2883138|T047|I82.549|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED TIBIAL VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED TIBIAL VEIN
C2883136|T047|I82.542|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF LEFT TIBIAL VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF LEFT TIBIAL VEIN
C2883137|T047|I82.543|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF TIBIAL VEIN, BILATERAL|CHRONIC EMBOLISM AND THROMBOSIS OF TIBIAL VEIN, BILATERAL
C2883135|T047|I82.541|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF RIGHT TIBIAL VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF RIGHT TIBIAL VEIN
C4267986|T047|E09.3529|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, UNSPECIFIED EYE|DRUG/CHEM DIAB W PROLIF DIAB RTNOP W TRCTN DTCH MACULA, UNSP
C2832557|T037|S06.812A|ICD10CM|INJURY OF RIGHT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|INJURY OF R INT CAROTID, INTCR W LOC OF 31-59 MIN, INIT
C2855944|T037|S68.129S|ICD10CM|PARTIAL TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF UNSPECIFIED FINGER, SEQUELA|PARTIAL TRAUMATIC MCP AMPUTATION OF UNSP FINGER, SEQUELA
C4267983|T047|E09.3521|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, RIGHT EYE|DRUG/CHEM DIAB W PROLIF DIAB RTNOP W TRCTN DTCH MACULA,R EYE
C4267985|T047|E09.3523|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, BILATERAL|DRUG/CHEM DIAB W PROLIF DIAB RTNOP W TRCTN DTCH MACULA, BI
C4267984|T047|E09.3522|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, LEFT EYE|DRUG/CHEM DIAB W PROLIF DIAB RTNOP W TRCTN DTCH MACULA,L EYE
C2905817|T037|X83.8XXA|ICD10CM|INTENTIONAL SELF-HARM BY OTHER SPECIFIED MEANS, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY OTHER SPECIFIED MEANS, INIT ENCNTR
C2858799|T037|S72.454A|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP SUPRCNDL FX W/O INTRCNDL EXTN LOWER END R FEMR, INIT
C2889097|T047|M02.861|ICD10CM|OTHER REACTIVE ARTHROPATHIES, RIGHT KNEE|OTHER REACTIVE ARTHROPATHIES, RIGHT KNEE
C2842049|T191|C49.8|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF CONNECTIVE AND SOFT TISSUE|PRIMARY MALIGNANT NEOPLASM OF TWO OR MORE CONTIGUOUS SITES OF CONNECTIVE AND SOFT TISSUE
C2889098|T047|M02.862|ICD10CM|OTHER REACTIVE ARTHROPATHIES, LEFT KNEE|OTHER REACTIVE ARTHROPATHIES, LEFT KNEE
C0348361|T191|C49.6|DMDICD10|MALIGNANT NEOPLASM OF CONNECTIVE AND SOFT TISSUE OF TRUNK, UNSPECIFIED|BOESARTIGE NEUBILDUNG: BINDEGEWEBE UND ANDERE WEICHTEILGEWEBE DES RUMPFES, NICHT NAEHER BEZEICHNET
C0864917|T191|C49.4|ICD10CM|MALIGNANT NEOPLASM OF CONNECTIVE AND SOFT TISSUE OF ABDOMEN|MALIGNANT NEOPLASM OF HYPOCHONDRIUM
C0864921|T191|C49.5|ICD10CM|MALIGNANT NEOPLASM OF CONNECTIVE AND SOFT TISSUE OF PELVIS|MALIGNANT NEOPLASM OF PERINEUM
C2889099|T047|M02.86|ICD10CM|OTHER REACTIVE ARTHROPATHIES, UNSPECIFIED KNEE|OTHER REACTIVE ARTHROPATHIES, KNEE
C3665405|T191|C49.3|ICD10CM|MALIGNANT NEOPLASM OF CONNECTIVE AND SOFT TISSUE OF THORAX|MALIGNANT NEOPLASM OF GREAT VESSELS
C2118406|T191||ICD10CM|MALIGNANT NEOPLASM OF CONNECTIVE AND SOFT TISSUE OF HEAD, FACE AND NECK
C2856724|T037|S72.033A|ICD10CM|DISPLACED MIDCERVICAL FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED MIDCERVICAL FRACTURE OF UNSP FEMUR, INIT
C2977161|T046|T87.1X9|ICD10CM|COMPLICATIONS OF REATTACHED (PART OF) UNSPECIFIED LOWER EXTREMITY|COMPLICATIONS OF REATTACHED (PART OF) UNSP LOWER EXTREMITY
C2856726|T037|S72.033C|ICD10CM|DISPLACED MIDCERVICAL FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL MIDCERVICAL FX UNSP FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2856725|T037|S72.033B|ICD10CM|DISPLACED MIDCERVICAL FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL MIDCERVICAL FX UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2858475|T037|S72.423B|ICD10CM|DISPLACED FRACTURE OF LATERAL CONDYLE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF LATERAL CONDYLE OF UNSP FEMR, 7THB
C2882410|T047|I63.539|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF UNSPECIFIED POSTERIOR CEREBRAL ARTERY|CEREB INFRC D/T UNSP OCCLS OR STENOS OF UNSP POST CEREB ART
C2843325|T037|S48.912A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT SHOULDER AND UPPER ARM, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|COMPLETE TRAUM AMP OF LEFT SHLDR/UP ARM, LEVEL UNSP, INIT
C2882409|T047|I63.532|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF LEFT POSTERIOR CEREBRAL ARTERY|CEREB INFRC D/T UNSP OCCLS OR STENOS OF LEFT POST CEREB ART
C4268491|T046|I63.533|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF BILATERAL POSTERIOR CEREBRAL ARTERIES|CEREB INFRC DUE TO UNSP OCCLS OR STENOS OF BI POST CEREB ART
C2882408|T047|I63.531|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF RIGHT POSTERIOR CEREBRAL ARTERY|CEREB INFRC D/T UNSP OCCLS OR STENOS OF RIGHT POST CEREB ART
C2884414|T037|T54.92XA|ICD10CM|TOXIC EFFECT OF UNSPECIFIED CORROSIVE SUBSTANCE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF UNSP CORROSIVE SUBSTANCE, SELF-HARM, INIT
C2889130|T047|M05.072|ICD10CM|FELTY'S SYNDROME, LEFT ANKLE AND FOOT|FELTY'S SYNDROME, LEFT ANKLE AND FOOT
C2889129|T047|M05.071|ICD10CM|FELTY'S SYNDROME, RIGHT ANKLE AND FOOT|FELTY'S SYNDROME, RIGHT ANKLE AND FOOT
C2889131|T047|M05.079|ICD10CM|FELTY'S SYNDROME, UNSPECIFIED ANKLE AND FOOT|FELTY'S SYNDROME, UNSPECIFIED ANKLE AND FOOT
C2843327|T037|S48.912S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT SHOULDER AND UPPER ARM, LEVEL UNSPECIFIED, SEQUELA|COMPLETE TRAUM AMP OF LEFT SHLDR/UP ARM, LEVEL UNSP, SEQUELA
C2858045|T037|S72.352A|ICD10CM|DISPLACED COMMINUTED FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED COMMINUTED FRACTURE OF SHAFT OF LEFT FEMUR, INIT
C2858047|T037|S72.352C|ICD10CM|DISPLACED COMMINUTED FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL COMMNT FX SHAFT OF L FEMR, INIT FOR OPN FX TYPE 3A/B/C
C2858046|T037|S72.352B|ICD10CM|DISPLACED COMMINUTED FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL COMMNT FX SHAFT OF L FEMUR, INIT FOR OPN FX TYPE I/2
C2884138|T037|T52.3X2S|ICD10CM|TOXIC EFFECT OF GLYCOLS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF GLYCOLS, INTENTIONAL SELF-HARM, SEQUELA
C2884544|T037|T56.5X2A|ICD10CM|TOXIC EFFECT OF ZINC AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF ZINC AND ITS COMPOUNDS, SELF-HARM, INIT
C2884136|T037|T52.3X2A|ICD10CM|TOXIC EFFECT OF GLYCOLS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF GLYCOLS, INTENTIONAL SELF-HARM, INIT ENCNTR
C2860127|T037|S79.102A|ICD10CM|UNSPECIFIED PHYSEAL FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP PHYSEAL FRACTURE OF LOWER END OF LEFT FEMUR, INIT
C2838151|T037|S32.443B|ICD10CM|DISPLACED FRACTURE OF POSTERIOR COLUMN [ILIOISCHIAL] OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISP FX OF POSTERIOR COLUMN OF UNSP ACETAB, INIT FOR OPN FX
C2838150|T037|S32.443A|ICD10CM|DISPLACED FRACTURE OF POSTERIOR COLUMN [ILIOISCHIAL] OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF POSTERIOR COLUMN OF UNSP ACETABULUM, INIT
C2884546|T037|T56.5X2S|ICD10CM|TOXIC EFFECT OF ZINC AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF ZINC AND ITS COMPOUNDS, SELF-HARM, SEQUELA
C2838358|T037|S32.492A|ICD10CM|OTHER SPECIFIED FRACTURE OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF LEFT ACETABULUM, INIT FOR CLOS FX
C2838359|T037|S32.492B|ICD10CM|OTHER SPECIFIED FRACTURE OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF LEFT ACETABULUM, INIT FOR OPN FX
C2890962|T037|T85.118A|ICD10CM|BREAKDOWN (MECHANICAL) OF OTHER IMPLANTED ELECTRONIC STIMULATOR OF NERVOUS SYSTEM, INITIAL ENCOUNTER|BRKDWN IMPLANTED ELECTRONIC STIMULATOR OF NERVOUS SYS, INIT
C2838616|T037|S34.101A|ICD10CM|UNSPECIFIED INJURY TO L1 LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY TO L1 LEVEL OF LUMBAR SPINAL CORD, INIT ENCNTR
C2876232|T037|T32.96|ICD10CM|CORROSIONS INVOLVING 90% OR MORE OF BODY SURFACE WITH 60-69% THIRD DEGREE CORROSION|CORROS 90%/MORE OF BODY SURFACE W 60-69% THIRD DEGREE CORROS
C2902137|T046|M87.835|ICD10CM|OTHER OSTEONECROSIS OF LEFT ULNA|OTHER OSTEONECROSIS OF LEFT ULNA
C2902136|T046|M87.834|ICD10CM|OTHER OSTEONECROSIS OF RIGHT ULNA|OTHER OSTEONECROSIS OF RIGHT ULNA
C2902139|T046|M87.837|ICD10CM|OTHER OSTEONECROSIS OF RIGHT CARPUS|OTHER OSTEONECROSIS OF RIGHT CARPUS
C2902138|T046|M87.836|ICD10CM|OTHER OSTEONECROSIS OF UNSPECIFIED ULNA|OTHER OSTEONECROSIS OF UNSPECIFIED ULNA
C2902133|T046|M87.831|ICD10CM|OTHER OSTEONECROSIS OF RIGHT RADIUS|OTHER OSTEONECROSIS OF RIGHT RADIUS
C2890891|T037|T84.69XA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL FIXATION DEVICE OF OTHER SITE, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INT FIX OF SITE, INIT
C2902135|T046|M87.833|ICD10CM|OTHER OSTEONECROSIS OF UNSPECIFIED RADIUS|OTHER OSTEONECROSIS OF UNSPECIFIED RADIUS
C2902134|T046|M87.832|ICD10CM|OTHER OSTEONECROSIS OF LEFT RADIUS|OTHER OSTEONECROSIS OF LEFT RADIUS
C4267849|T191|C81.26|ICD10CM|MIXED CELLULARITY HODGKIN LYMPHOMA, INTRAPELVIC LYMPH NODES|MIXED CELLULARITY HODGKIN LYMPHOMA, INTRAPELVIC LYMPH NODES
C2902141|T046|M87.839|ICD10CM|OTHER OSTEONECROSIS OF UNSPECIFIED CARPUS|OTHER OSTEONECROSIS OF UNSPECIFIED CARPUS
C2902140|T046|M87.838|ICD10CM|OTHER OSTEONECROSIS OF LEFT CARPUS|OTHER OSTEONECROSIS OF LEFT CARPUS
C2858678|T037|S72.443A|ICD10CM|DISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF LOWER EPIPHYSIS (SEPARATION) OF UNSP FEMUR, INIT
C2889323|T047|M05.672|ICD10CM|RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF LEFT ANK/FT W INVOLV OF ORGANS AND SYSTEMS
C0477367|T047|G36.8|DMDICD10|OTHER SPECIFIED ACUTE DISSEMINATED DEMYELINATION|SONSTIGE NAEHER BEZEICHNETE AKUTE DISSEMINIERTE DEMYELINISATION
C0477368|T047|G36.9|DMDICD10|ACUTE DISSEMINATED DEMYELINATION, UNSPECIFIED|AKUTE DISSEMINIERTE DEMYELINISATION, NICHT NAEHER BEZEICHNET
C2891322|T037|T87.1X2|ICD10CM|COMPLICATIONS OF REATTACHED (PART OF) LEFT LOWER EXTREMITY|COMPLICATIONS OF REATTACHED (PART OF) LEFT LOWER EXTREMITY
C1395170|T047||ICD10CM|NEUROMYELITIS OPTICA [DEVIC]
C0349367|T047|G36.1|DMDICD10|ACUTE AND SUBACUTE HEMORRHAGIC LEUKOENCEPHALITIS [HURST]|AKUTE UND SUBAKUTE HAEMORRHAGISCHE LEUKOENZEPHALITIS [HURST]
C2857068|T037|S72.092A|ICD10CM|OTHER FRACTURE OF HEAD AND NECK OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF HEAD AND NECK OF LEFT FEMUR, INIT
C2857069|T037|S72.092B|ICD10CM|OTHER FRACTURE OF HEAD AND NECK OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|OTH FX HEAD/NECK OF LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C2857070|T037|S72.092C|ICD10CM|OTHER FRACTURE OF HEAD AND NECK OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|OTH FX HEAD/NECK OF LEFT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2874296|T047|E80.3|ICD10CM|DEFECTS OF CATALASE AND PEROXIDASE|ACATALASIA [TAKAHARA]
C0260976|T037|E801|ICD9CM|PORPHYRIA CUTANEA TARDA|RAILWAY ACCIDENT INVOLVING COLLISION WITH OTHER OBJECT
C0260969|T037|E800|ICD9CM|HEREDITARY ERYTHROPOIETIC PORPHYRIA|RAILWAY ACCIDENT INVOLVING COLLISION WITH ROLLING STOCK
C2882187|T047|I25.729|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS ARTERY CORONARY ARTERY BYPASS GRAFT(S) WITH UNSPECIFIED ANGINA PECTORIS|ATHSCL AUTOLOGOUS ARTERY CABG W UNSP ANGINA PECTORIS
C2882186|T047|I25.728|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS ARTERY CORONARY ARTERY BYPASS GRAFT(S) WITH OTHER FORMS OF ANGINA PECTORIS|ATHSCL AUTOLOGOUS ARTERY CABG W OTH ANGINA PECTORIS
C2837996|T191|C43.59|ICD10CM|MALIGNANT MELANOMA OF OTHER PART OF TRUNK|MALIGNANT MELANOMA OF OTHER PART OF TRUNK
C0348426|T191|D32|DMDICD10|BENIGN NEOPLASM OF MENINGES, UNSPECIFIED|GUTARTIGE NEUBILDUNG DER MENINGEN
C2882184|T047|I25.720|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS ARTERY CORONARY ARTERY BYPASS GRAFT(S) WITH UNSTABLE ANGINA PECTORIS|ATHSCL AUTOLOGOUS ARTERY CABG W UNSTABLE ANGINA PECTORIS
C0684503|T191|C43.52|ICD10CM|MALIGNANT MELANOMA OF SKIN OF BREAST|MALIGNANT MELANOMA OF SKIN OF BREAST
C2837995|T191|C43.51|ICD10CM|MALIGNANT MELANOMA OF ANAL SKIN|MALIGNANT MELANOMA OF ANAL SKIN
C4267926|T047|E08.3521|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, RIGHT EYE|DIAB WITH PROLIF DIAB RTNOP WITH TRCTN DTCH MACULA, R EYE
C4267927|T047|E08.3522|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, LEFT EYE|DIAB WITH PROLIF DIAB RTNOP WITH TRCTN DTCH MACULA, LEFT EYE
C4267928|T047|E08.3523|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, BILATERAL|DIAB WITH PROLIF DIABETIC RTNOP WITH TRCTN DTCH MACULA, BI
C2877046|T037|T38.2X2A|ICD10CM|POISONING BY ANTITHYROID DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ANTITHYROID DRUGS, INTENTIONAL SELF-HARM, INIT
C4267929|T047|E08.3529|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT INVOLVING THE MACULA, UNSPECIFIED EYE|DIAB WITH PROLIF DIABETIC RTNOP WITH TRCTN DTCH MACULA, UNSP
C2853978|T191|C84.68|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-POSITIVE, LYMPH NODES OF MULTIPLE SITES|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-POS, NODES MULT SITE
C2853979|T191|C84.69|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-POSITIVE, EXTRANODAL AND SOLID ORGAN SITES|ANAPLSTC LG CELL LYMPH, ALK-POS, EXTRNOD AND SOLID ORG SITES
C2853974|T191|C84.64|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-POSITIVE, LYMPH NODES OF AXILLA AND UPPER LIMB|ANAPLSTC LG CELL LYMPH, ALK-POS, NODES OF AXLA AND UPR LIMB
C2853975|T191|C84.65|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-POSITIVE, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|ANAPLSTC LG CELL LYMPH, ALK-POS, NODES OF ING RGN & LOW LMB
C2853976|T191|C84.66|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-POSITIVE, INTRAPELVIC LYMPH NODES|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-POS, INTRAPELV NODES
C2853977|T191||ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-POSITIVE, SPLEEN
C2853970|T191|C84.60|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-POSITIVE, UNSPECIFIED SITE|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-POSITIVE, UNSP SITE
C2853971|T191|C84.61|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-POSITIVE, LYMPH NODES OF HEAD, FACE, AND NECK|ANAPLSTC LG CELL LYMPH, ALK-POS, NODES OF HEAD, FACE, AND NK
C2853972|T191|C84.62|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-POSITIVE, INTRATHORACIC LYMPH NODES|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-POS, INTRATHORAC NODES
C2853973|T191|C84.63|ICD10CM|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-POSITIVE, INTRA-ABDOMINAL LYMPH NODES|ANAPLASTIC LARGE CELL LYMPHOMA, ALK-POS, INTRA-ABD NODES
C4268144|T047|E13.3419|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|OTH DIABETES WITH SEVERE NONP RTNOP WITH MACULAR EDEMA, UNSP
C2861587|T191|C92.21|ICD10CM|ATYPICAL CHRONIC MYELOID LEUKEMIA, BCR/ABL-NEGATIVE, IN REMISSION|ATYPICAL CHRONIC MYELOID LEUKEMIA, BCR/ABL-NEG, IN REMISSION
C4268141|T047|E13.3411|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|OTH DIAB WITH SEVERE NONP RTNOP WITH MACULAR EDEMA, R EYE
C4268142|T047|E13.3412|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|OTH DIAB WITH SEVERE NONP RTNOP WITH MACULAR EDEMA, LEFT EYE
C4268143|T047|E13.3413|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|OTH DIABETES WITH SEVERE NONP RTNOP WITH MACULAR EDEMA, BI
C2890463|T037|T84.032A|ICD10CM|MECHANICAL LOOSENING OF INTERNAL RIGHT KNEE PROSTHETIC JOINT, INITIAL ENCOUNTER|MECH LOOSENING OF INTERNAL RIGHT KNEE PROSTHETIC JOINT, INIT
C3264362|T047|A41.01|ICD10CM|SEPSIS DUE TO METHICILLIN SUSCEPTIBLE STAPHYLOCOCCUS AUREUS|SEPSIS DUE TO METHICILLIN SUSCEPTIBLE STAPHYLOCOCCUS AUREUS
C3164390|T047||ICD10CM|SEPSIS DUE TO METHICILLIN RESISTANT STAPHYLOCOCCUS AUREUS
C2882818|T047|I70.428|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, OTHER EXTREMITY|ATHSCL AUTOL VEIN BYPASS OF THE EXTRM W REST PAIN, OTH EXTRM
C2882819|T047|I70.429|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, UNSPECIFIED EXTREMITY|ATHSCL AUTOL VEIN BYPASS OF EXTRM W REST PAIN, UNSP EXTRM
C2882815|T047|I70.421|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, RIGHT LEG|ATHSCL AUTOL VEIN BYPASS OF THE EXTRM W REST PAIN, RIGHT LEG
C2882816|T047|I70.422|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, LEFT LEG|ATHSCL AUTOL VEIN BYPASS OF THE EXTRM W REST PAIN, LEFT LEG
C2882817|T047|I70.423|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, BILATERAL LEGS|ATHSCL AUTOL VEIN BYPASS OF THE EXTRM W REST PAIN, BI LEGS
C2832018|T037|S06.2X1S|ICD10CM|DIFFUSE TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|DIFFUSE TBI W LOC OF 30 MINUTES OR LESS, SEQUELA
C0276308|T047|B06.82|ICD10CM|RUBELLA ARTHRITIS|RUBELLA ARTHRITIS
C2877664|T037|T40.4X2S|ICD10CM|POISONING BY OTHER SYNTHETIC NARCOTICS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH SYNTHETIC NARCOTICS, SELF-HARM, SEQUELA
C2833256|T037|S12.121A|ICD10CM|OTHER NONDISPLACED DENS FRACTURE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH NONDISPLACED DENS FRACTURE, INIT FOR CLOS FX
C2835845|T037|S24.152A|ICD10CM|OTHER INCOMPLETE LESION AT T2-T6 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|OTH INCOMPLETE LESION AT T2-T6, INIT
C2835846|T037|S24.152D|ICD10CM|OTHER INCOMPLETE LESION AT T2-T6 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|OTH INCOMPLETE LESION AT T2-T6, SUBS
C0264797|T047|B33.24|ICD10CM|VIRAL CARDIOMYOPATHY|VIRAL CARDIOMYOPATHY
C2877662|T037|T40.4X2A|ICD10CM|POISONING BY OTHER SYNTHETIC NARCOTICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH SYNTHETIC NARCOTICS, SELF-HARM, INIT
C0494266|T047|D84.8|DMDICD10|OTHER SPECIFIED IMMUNODEFICIENCIES|SONSTIGE NAEHER BEZEICHNETE IMMUNDEFEKTE
C2876132|T037|T31.22|ICD10CM|BURNS INVOLVING 20-29% OF BODY SURFACE WITH 20-29% THIRD DEGREE BURNS|BURNS OF 20-29% OF BODY SURFACE W 20-29% THIRD DEGREE BURNS
C2838473|T037|S32.691B|ICD10CM|OTHER SPECIFIED FRACTURE OF RIGHT ISCHIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF RIGHT ISCHIUM, INIT ENCNTR FOR OPEN FRACTURE
C2838472|T037|S32.691A|ICD10CM|OTHER SPECIFIED FRACTURE OF RIGHT ISCHIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF RIGHT ISCHIUM, INIT FOR CLOS FX
C2838072|T037|S32.424B|ICD10CM|NONDISPLACED FRACTURE OF POSTERIOR WALL OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP FX OF POST WALL OF RIGHT ACETAB, INIT FOR OPN FX
C2832389|T037|S06.380S|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF BRAINSTEM WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|CONTUS/LAC/HEM BRAINSTEM W/O LOSS OF CONSCIOUSNESS, SEQUELA
C2901817|T047|M86.172|ICD10CM|OTHER ACUTE OSTEOMYELITIS, LEFT ANKLE AND FOOT|OTHER ACUTE OSTEOMYELITIS, LEFT ANKLE AND FOOT
C0036337|T048|F25|DMDICD10|SCHIZOAFFECTIVE DISORDER, UNSPECIFIED|SCHIZOAFFEKTIVE STOERUNGEN
C0349201|T048|F25.8|DMDICD10|OTHER SCHIZOAFFECTIVE DISORDERS|SONSTIGE SCHIZOAFFEKTIVE STOERUNGEN
C4269529|T037|S02.650S|ICD10CM|FRACTURE OF ANGLE OF MANDIBLE, UNSPECIFIED SIDE, SEQUELA|FRACTURE OF ANGLE OF MANDIBLE, UNSPECIFIED SIDE, SEQUELA
C1405641|T048||ICD10CM|SCHIZOAFFECTIVE DISORDER, DEPRESSIVE TYPE
C2874858|T048|F25.0|ICD10CM|SCHIZOAFFECTIVE DISORDER, BIPOLAR TYPE|SCHIZOAFFECTIVE PSYCHOSIS, BIPOLAR TYPE
C2832387|T037|S06.380A|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF BRAINSTEM WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|CONTUS/LAC/HEM BRAINSTEM W/O LOSS OF CONSCIOUSNESS, INIT
C4269524|T037|S02.650A|ICD10CM|FRACTURE OF ANGLE OF MANDIBLE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF ANGLE OF MANDIBLE, UNSPECIFIED SIDE, INIT
C4269525|T037|S02.650B|ICD10CM|FRACTURE OF ANGLE OF MANDIBLE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF ANGLE OF MANDIBLE, UNSPECIFIED SIDE, 7THB
C2878765|T037|T44.1X2S|ICD10CM|POISONING BY OTHER PARASYMPATHOMIMETICS [CHOLINERGICS], INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH PARASYMPATHOMIMETICS, SELF-HARM, SEQUELA
C2885801|T037|T63.632S|ICD10CM|TOXIC EFFECT OF CONTACT WITH SEA ANEMONE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CONTACT W SEA ANEMONE, SELF-HARM, SEQUELA
C4236944|T048|F10.97|ICD10CM|ALCOHOL USE, UNSPECIFIED WITH ALCOHOL-INDUCED PERSISTING DEMENTIA|ALCOHOL-INDUCED MAJOR NEUROCOGNITIVE DISORDER, NONAMNESTIC-CONFABULATORY TYPE, WITHOUT USE DISORDER
C2889268|T047|M05.519|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER|RHEU POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP SHOULDER
C4268214|T048|F10.94|ICD10CM|ALCOHOL USE, UNSPECIFIED WITH ALCOHOL-INDUCED MOOD DISORDER|ALCOHOL INDUCED BIPOLAR OR RELATED DISORDER, WITHOUT USE DISORDER
C2885748|T037|T63.592S|ICD10CM|TOXIC EFFECT OF CONTACT WITH OTHER VENOMOUS FISH, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CONTACT W OTH VENOM FISH, SLF-HRM, SEQUELA
C2874420|T048|F10.99|ICD10CM|ALCOHOL USE, UNSPECIFIED WITH UNSPECIFIED ALCOHOL-INDUCED DISORDER|ALCOHOL USE, UNSP WITH UNSPECIFIED ALCOHOL-INDUCED DISORDER
C2889266|T047|M05.511|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT SHOULDER|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF R SHOULDER
C2889267|T047|M05.512|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT SHOULDER|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF L SHOULDER
C2885799|T037|T63.632A|ICD10CM|TOXIC EFFECT OF CONTACT WITH SEA ANEMONE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CONTACT W SEA ANEMONE, SELF-HARM, INIT
C2878763|T037|T44.1X2A|ICD10CM|POISONING BY OTHER PARASYMPATHOMIMETICS [CHOLINERGICS], INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH PARASYMPATHOMIMETICS, SELF-HARM, INIT
C2889637|T047|M08.939|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, UNSPECIFIED WRIST|JUVENILE ARTHRITIS, UNSPECIFIED, UNSPECIFIED WRIST
C2885746|T037|T63.592A|ICD10CM|TOXIC EFFECT OF CONTACT WITH OTHER VENOMOUS FISH, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CONTACT W OTH VENOMOUS FISH, SELF-HARM, INIT
C2889635|T047|M08.931|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, RIGHT WRIST|JUVENILE ARTHRITIS, UNSPECIFIED, RIGHT WRIST
C2889636|T047|M08.932|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, LEFT WRIST|JUVENILE ARTHRITIS, UNSPECIFIED, LEFT WRIST
C2878791|T037|T44.2X2S|ICD10CM|POISONING BY GANGLIONIC BLOCKING DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY GANGLIONIC BLOCKING DRUGS, SELF-HARM, SEQUELA
C2874479|T048|F12.159|ICD10CM|CANNABIS ABUSE WITH PSYCHOTIC DISORDER, UNSPECIFIED|CANNABIS ABUSE WITH PSYCHOTIC DISORDER, UNSPECIFIED
C2874284|T047|E76.29|ICD10CM|OTHER MUCOPOLYSACCHARIDOSES|MUCOPOLYSACCHARIDOSIS, TYPES VI, VII
C2874254|T047|E71.53|ICD10CM|OTHER GROUP 2 PEROXISOMAL DISORDERS|OTHER GROUP 2 PEROXISOMAL DISORDERS
C2874282|T047|E76.22|ICD10CM|SANFILIPPO MUCOPOLYSACCHARIDOSES|SANFILIPPO MUCOPOLYSACCHARIDOSES
C4268105|T047|E11.3539|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, UNSPECIFIED EYE|TYPE 2 DIAB W PROLIF DIAB RTNOP WITH TRCTN DTCH N-MCLA, UNSP
C2878789|T037|T44.2X2A|ICD10CM|POISONING BY GANGLIONIC BLOCKING DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY GANGLIONIC BLOCKING DRUGS, SELF-HARM, INIT
C2832676|T037|S06.9X1A|ICD10CM|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|UNSP INTRACRANIAL INJURY W LOC OF 30 MINUTES OR LESS, INIT
C2977942|T191|C65.2|ICD10CM|MALIGNANT NEOPLASM OF LEFT RENAL PELVIS|MALIGNANT NEOPLASM OF LEFT RENAL PELVIS
C4268102|T047|E11.3531|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, RIGHT EYE|TYPE 2 DIAB W PROLIF DIAB RTNOP W TRCTN DTCH N-MCLA, R EYE
C2832072|T037|S06.304S|ICD10CM|UNSPECIFIED FOCAL TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, SEQUELA|UNSP FOCAL TBI W LOC OF 6 HOURS TO 24 HOURS, SEQUELA
C4268104|T047|E11.3533|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, BILATERAL|TYPE 2 DIAB W PROLIF DIAB RTNOP WITH TRCTN DTCH N-MCLA, BI
C4268103|T047|E11.3532|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, LEFT EYE|TYPE 2 DIAB W PROLIF DIAB RTNOP W TRCTN DTCH N-MCLA, L EYE
C2838171|T037|S32.446A|ICD10CM|NONDISPLACED FRACTURE OF POSTERIOR COLUMN [ILIOISCHIAL] OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF POSTERIOR COLUMN OF UNSP ACETABULUM, INIT
C2858576|T037|S72.433A|ICD10CM|DISPLACED FRACTURE OF MEDIAL CONDYLE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF MEDIAL CONDYLE OF UNSP FEMUR, INIT FOR CLOS FX
C2858578|T037|S72.433C|ICD10CM|DISPLACED FRACTURE OF MEDIAL CONDYLE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF MED CONDYLE OF UNSP FEMR, 7THC
C2858577|T037|S72.433B|ICD10CM|DISPLACED FRACTURE OF MEDIAL CONDYLE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF MED CONDYLE OF UNSP FEMR, 7THB
C2837653|T037|S32.059A|ICD10CM|UNSPECIFIED FRACTURE OF FIFTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF FIFTH LUMBAR VERTEBRA, INIT FOR CLOS FX
C2837654|T037|S32.059B|ICD10CM|UNSPECIFIED FRACTURE OF FIFTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF FIFTH LUMBAR VERTEBRA, INIT FOR OPN FX
C4268015|T047|E10.3291|ICD10CM|TYPE 1 DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|TYPE 1 DIAB WITH MILD NONP RTNOP WITHOUT MCLR EDEMA, R EYE
C2874946|T048|F40.248|ICD10CM|OTHER SITUATIONAL TYPE PHOBIA|OTHER SITUATIONAL TYPE PHOBIA
C4268016|T047|E10.3292|ICD10CM|TYPE 1 DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|TYPE 1 DIAB WITH MILD NONP RTNOP WITHOUT MCLR EDEMA, L EYE
C2905786|T037|X81.8XXA|ICD10CM|INTENTIONAL SELF-HARM BY JUMPING OR LYING IN FRONT OF OTHER MOVING OBJECT, INITIAL ENCOUNTER|SLF-HRM BY JUMPING OR LYING IN FRONT OF MOVING OBJECT, INIT
C0348499|T047|E85.8|DMDICD10|OTHER AMYLOIDOSIS|SONSTIGE AMYLOIDOSE
C2874945|T048|F40.242|ICD10CM|FEAR OF BRIDGES|FEAR OF BRIDGES
C0424184|T048|F40.243|ICD10CM|FEAR OF FLYING|FEAR OF FLYING
C0008909|T048|F40.240|ICD10CM|CLAUSTROPHOBIA|CLAUSTROPHOBIA
C0233701|T048|F40.241|ICD10CM|ACROPHOBIA|ACROPHOBIA
C2205119|T191||ICD10CM|MALIGNANT CARCINOID TUMOR OF THE RECTUM
C2349319|T191||ICD10CM|MALIGNANT CARCINOID TUMOR OF THE CECUM
C2901887|T047|M86.471|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, RIGHT ANKLE AND FOOT|CHRONIC OSTEOMYELITIS W DRAINING SINUS, RIGHT ANKLE AND FOOT
C2062529|T191||ICD10CM|MALIGNANT CARCINOID TUMOR OF THE APPENDIX
C2883031|T047|I71.9|ICD10CM|AORTIC ANEURYSM OF UNSPECIFIED SITE, WITHOUT RUPTURE|AORTIC ANEURYSM OF UNSPECIFIED SITE, WITHOUT RUPTURE
C0741160|T047|I71.8|DMDICD10|AORTIC ANEURYSM OF UNSPECIFIED SITE, RUPTURED|AORTENANEURYSMA NICHT NAEHER BEZEICHNETER LOKALISATION, RUPTURIERT
C0496947|T191|D44.6|DMDICD10|NEOPLASM OF UNCERTAIN BEHAVIOR OF CAROTID BODY|NEUBILDUNG UNSICHEREN ODER UNBEKANNTEN VERHALTENS: GLOMUS CAROTICUM
C0265012|T047|I71.3|DMDICD10|ABDOMINAL AORTIC ANEURYSM, RUPTURED|ANEURYSMA DER AORTA ABDOMINALIS, RUPTURIERT
C3251816|T020|I71.2|DMDICD10|THORACIC AORTIC ANEURYSM, WITHOUT RUPTURE|ANEURYSMA DER AORTA THORACICA, OHNE ANGABE EINER RUPTUR
C0265010|T047|I71.1|DMDICD10|THORACIC AORTIC ANEURYSM, RUPTURED|ANEURYSMA DER AORTA THORACICA, RUPTURIERT
C2873710|T191|D44.7|ICD10CM|NEOPLASM OF UNCERTAIN BEHAVIOR OF AORTIC BODY AND OTHER PARAGANGLIA|NEOPLASM OF UNCRT BEHAV OF AORTIC BODY AND OTH PARAGANGLIA
C2883030|T047|I71.6|ICD10CM|THORACOABDOMINAL AORTIC ANEURYSM, WITHOUT RUPTURE|THORACOABDOMINAL AORTIC ANEURYSM, WITHOUT RUPTURE
C1305122|T047|I71.5|DMDICD10|THORACOABDOMINAL AORTIC ANEURYSM, RUPTURED|AORTENANEURYSMA, THORAKOABDOMINAL, RUPTURIERT
C0265011|T020|I71.4|DMDICD10|ABDOMINAL AORTIC ANEURYSM, WITHOUT RUPTURE|ANEURYSMA DER AORTA ABDOMINALIS, OHNE ANGABE EINER RUPTUR
C2884978|T037|T59.892A|ICD10CM|TOXIC EFFECT OF OTHER SPECIFIED GASES, FUMES AND VAPORS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF GASES, FUMES AND VAPORS, SELF-HARM, INIT
C2859097|T037|S72.91XB|ICD10CM|UNSPECIFIED FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP FRACTURE OF RIGHT FEMUR, INIT FOR OPN FX TYPE I/2
C2834027|T037|S14.149S|ICD10CM|BROWN-SEQUARD SYNDROME AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, SEQUELA|BROWN-SEQUARD SYND AT UNSP LEVEL OF CERV SPINAL CORD, SQLA
C2902095|T046|M87.338|ICD10CM|OTHER SECONDARY OSTEONECROSIS OF LEFT CARPUS|OTHER SECONDARY OSTEONECROSIS OF LEFT CARPUS
C2902096|T046|M87.339|ICD10CM|OTHER SECONDARY OSTEONECROSIS OF UNSPECIFIED CARPUS|OTHER SECONDARY OSTEONECROSIS OF UNSPECIFIED CARPUS
C2832070|T037|S06.304A|ICD10CM|UNSPECIFIED FOCAL TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|UNSP FOCAL TBI W LOC OF 6 HOURS TO 24 HOURS, INIT
C2902089|T046|M87.332|ICD10CM|OTHER SECONDARY OSTEONECROSIS OF LEFT RADIUS|OTHER SECONDARY OSTEONECROSIS OF LEFT RADIUS
C2902090|T046|M87.333|ICD10CM|OTHER SECONDARY OSTEONECROSIS OF UNSPECIFIED RADIUS|OTHER SECONDARY OSTEONECROSIS OF UNSPECIFIED RADIUS
C4270227|T046|T83.038A|ICD10CM|LEAKAGE OF OTHER URINARY CATHETER, INITIAL ENCOUNTER|LEAKAGE OF OTHER URINARY CATHETER, INITIAL ENCOUNTER
C2902088|T046|M87.331|ICD10CM|OTHER SECONDARY OSTEONECROSIS OF RIGHT RADIUS|OTHER SECONDARY OSTEONECROSIS OF RIGHT RADIUS
C2902093|T046|M87.336|ICD10CM|OTHER SECONDARY OSTEONECROSIS OF UNSPECIFIED ULNA|OTHER SECONDARY OSTEONECROSIS OF UNSPECIFIED ULNA
C2902094|T046|M87.337|ICD10CM|OTHER SECONDARY OSTEONECROSIS OF RIGHT CARPUS|OTHER SECONDARY OSTEONECROSIS OF RIGHT CARPUS
C2902091|T046|M87.334|ICD10CM|OTHER SECONDARY OSTEONECROSIS OF RIGHT ULNA|OTHER SECONDARY OSTEONECROSIS OF RIGHT ULNA
C2902092|T046|M87.335|ICD10CM|OTHER SECONDARY OSTEONECROSIS OF LEFT ULNA|OTHER SECONDARY OSTEONECROSIS OF LEFT ULNA
C2835219|T037|S22.019B|ICD10CM|UNSPECIFIED FRACTURE OF FIRST THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF FIRST THORACIC VERTEBRA, INIT FOR OPN FX
C2835218|T037|S22.019A|ICD10CM|UNSPECIFIED FRACTURE OF FIRST THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF FIRST THORACIC VERTEBRA, INIT FOR CLOS FX
C2833649|T037|S12.8XXA|ICD10CM|FRACTURE OF OTHER PARTS OF NECK, INITIAL ENCOUNTER|FRACTURE OF OTHER PARTS OF NECK, INITIAL ENCOUNTER
C2883039|T046|I74.10|ICD10CM|EMBOLISM AND THROMBOSIS OF UNSPECIFIED PARTS OF AORTA|EMBOLISM AND THROMBOSIS OF UNSPECIFIED PARTS OF AORTA
C0155750|T046||ICD10CM|EMBOLISM AND THROMBOSIS OF THORACIC AORTA
C2832215|T037|S06.339A|ICD10CM|CONTUSION AND LACERATION OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|CONTUS/LAC CEREB, W LOC OF UNSP DURATION, INIT
C2882705|T047|I70.222|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES WITH REST PAIN, LEFT LEG|ATHSCL NATIVE ARTERIES OF EXTREMITIES W REST PAIN, LEFT LEG
C2882706|T047|I70.223|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES WITH REST PAIN, BILATERAL LEGS|ATHSCL NATIVE ARTERIES OF EXTRM W REST PAIN, BILATERAL LEGS
C2883040|T046|I74.19|ICD10CM|EMBOLISM AND THROMBOSIS OF OTHER PARTS OF AORTA|EMBOLISM AND THROMBOSIS OF OTHER PARTS OF AORTA
C2857823|T037|S72.331B|ICD10CM|DISPLACED OBLIQUE FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL OBLIQUE FX SHAFT OF R FEMUR, INIT FOR OPN FX TYPE I/2
C2857824|T037|S72.331C|ICD10CM|DISPLACED OBLIQUE FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL OBLIQUE FX SHAFT OF R FEMR, 7THC
C2857822|T037|S72.331A|ICD10CM|DISPLACED OBLIQUE FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED OBLIQUE FRACTURE OF SHAFT OF RIGHT FEMUR, INIT
C2879696|T037|T47.1X2A|ICD10CM|POISONING BY OTHER ANTACIDS AND ANTI-GASTRIC-SECRETION DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY OTH ANTACIDS & ANTI-GSTRC-SEC DRUGS, SLF-HRM, INIT
C2874058|T047|E10.618|ICD10CM|TYPE 1 DIABETES MELLITUS WITH OTHER DIABETIC ARTHROPATHY|TYPE 1 DIABETES MELLITUS WITH OTHER DIABETIC ARTHROPATHY
C2858183|T037|S72.364B|ICD10CM|NONDISPLACED SEGMENTAL FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP SEG FX SHAFT OF R FEMUR, INIT FOR OPN FX TYPE I/2
C2858184|T037|S72.364C|ICD10CM|NONDISPLACED SEGMENTAL FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP SEG FX SHAFT OF R FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C4268667|T046|K90.49|ICD10CM|MALABSORPTION DUE TO INTOLERANCE, NOT ELSEWHERE CLASSIFIED|MALABSORPTION DUE TO INTOLERANCE TO STARCH
C2896633|T046|M80.079A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, UNSPECIFIED ANKLE AND FOOT, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, UNSP ANK/FT, INIT
C2874057|T047|E10.610|ICD10CM|TYPE 1 DIABETES MELLITUS WITH DIABETIC NEUROPATHIC ARTHROPATHY|TYPE 1 DIABETES MELLITUS W DIABETIC NEUROPATHIC ARTHROPATHY
C2879698|T037|T47.1X2S|ICD10CM|POISONING BY OTHER ANTACIDS AND ANTI-GASTRIC-SECRETION DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY OTH ANTACIDS & ANTI-GSTRC-SEC DRUGS, SLF-HRM, SQLA
C2857224|T037|S72.115C|ICD10CM|NONDISPLACED FRACTURE OF GREATER TROCHANTER OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF GREATER TROCHANTER OF L FEMR, 7THC
C2838694|T037|S34.131D|ICD10CM|COMPLETE LESION OF SACRAL SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION OF SACRAL SPINAL CORD, SUBSEQUENT ENCOUNTER
C2838693|T037|S34.131A|ICD10CM|COMPLETE LESION OF SACRAL SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION OF SACRAL SPINAL CORD, INITIAL ENCOUNTER
C2890712|T037|T84.220A|ICD10CM|DISPLACEMENT OF INTERNAL FIXATION DEVICE OF BONES OF HAND AND FINGERS, INITIAL ENCOUNTER|DISPLACEMENT OF INT FIX OF BONES OF HAND AND FINGERS, INIT
C2838695|T037|S34.131S|ICD10CM|COMPLETE LESION OF SACRAL SPINAL CORD, SEQUELA|COMPLETE LESION OF SACRAL SPINAL CORD, SEQUELA
C2900982|T046|M84.446A|ICD10CM|PATHOLOGICAL FRACTURE, UNSPECIFIED FINGER(S), INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, UNSP FINGER(S), INIT FOR FX
C0342174|T047|E06.0|ICD10CM|ACUTE THYROIDITIS|ABSCESS OF THYROID
C2848454|T037|S58.921A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT FOREARM, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF R FOREARM, LEVEL UNSP, INIT
C2848456|T037|S58.921S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT FOREARM, LEVEL UNSPECIFIED, SEQUELA|PARTIAL TRAUMATIC AMP OF R FOREARM, LEVEL UNSP, SEQUELA
C0153470|T191|C26.1|DMDICD10|MALIGNANT NEOPLASM OF SPLEEN|BOESARTIGE NEUBILDUNG: MILZ
C0346627|T191|C26.0|DMDICD10|MALIGNANT NEOPLASM OF INTESTINAL TRACT, PART UNSPECIFIED|BOESARTIGE NEUBILDUNG: INTESTINALTRAKT, TEIL NICHT NAEHER BEZEICHNET
C2889054|T047|M02.322|ICD10CM|REITER'S DISEASE, LEFT ELBOW|REITER'S DISEASE, LEFT ELBOW
C2889053|T047|M02.321|ICD10CM|REITER'S DISEASE, RIGHT ELBOW|REITER'S DISEASE, RIGHT ELBOW
C0864885|T191|C26.9|ICD10CM|MALIGNANT NEOPLASM OF ILL-DEFINED SITES WITHIN THE DIGESTIVE SYSTEM|MALIGNANT NEOPLASM OF ALIMENTARY CANAL OR TRACT NOS
C2860164|T037|S79.121A|ICD10CM|SALTER-HARRIS TYPE II PHYSEAL FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SLTR-HARIS TYPE II PHYSEAL FX LOWER END OF RIGHT FEMUR, INIT
C2889055|T047|M02.329|ICD10CM|REITER'S DISEASE, UNSPECIFIED ELBOW|REITER'S DISEASE, UNSPECIFIED ELBOW
C2888392|T047|L89.219|ICD10CM|PRESSURE ULCER OF RIGHT HIP, UNSPECIFIED STAGE|PRESSURE ULCER OF RIGHT HIP, UNSPECIFIED STAGE
C2888389|T047|L89.214|ICD10CM|PRESSURE ULCER OF RIGHT HIP, STAGE 4|PRESSURE ULCER OF RIGHT HIP, STAGE 4
C2888377|T047||ICD10CM|PRESSURE ULCER OF RIGHT HIP, UNSTAGEABLE
C2888380|T047|L89.211|ICD10CM|PRESSURE ULCER OF RIGHT HIP, STAGE 1|PRESSURE ULCER OF RIGHT HIP, STAGE 1
C2888383|T047|L89.212|ICD10CM|PRESSURE ULCER OF RIGHT HIP, STAGE 2|PRESSURE ULCER OF RIGHT HIP, STAGE 2
C2888386|T047|L89.213|ICD10CM|PRESSURE ULCER OF RIGHT HIP, STAGE 3|PRESSURE ULCER OF RIGHT HIP, STAGE 3
C2874215|T047|E42|ICD10CM|MARASMIC KWASHIORKOR|SEVERE PROTEIN-CALORIE MALNUTRITION WITH SIGNS OF BOTH KWASHIORKOR AND MARASMUS
C2874216|T047|E43|ICD10CM|UNSPECIFIED SEVERE PROTEIN-CALORIE MALNUTRITION|UNSPECIFIED SEVERE PROTEIN-CALORIE MALNUTRITION
C0022806|T047|E40|DMDICD10|KWASHIORKOR|KWASHIORKOR
C0086588|T047|E41|DMDICD10|NUTRITIONAL MARASMUS|ALIMENTAERER MARASMUS
C2875092|T047|G40.201|ICD10CM|LOCALIZATION-RELATED (FOCAL) (PARTIAL) SYMPTOMATIC EPILEPSY AND EPILEPTIC SYNDROMES WITH COMPLEX PARTIAL SEIZURES, NOT INTRACTABLE, WITH STATUS EPILEPTICUS|LOCAL-REL SYMPTC EPI W CMPLX PRT SEIZ, NOT NTRCT, W STAT EPI
C2874220|T047|E45|ICD10CM|RETARDED DEVELOPMENT FOLLOWING PROTEIN-CALORIE MALNUTRITION|RETARDED DEVELOPMENT FOLLOWING PROTEIN-CALORIE MALNUTRITION
C2887923|T047||ICD10CM|TOXIC LIVER DISEASE WITH HEPATIC NECROSIS, WITH COMA
C2889238|T047|M05.422|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT ELBOW|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2890575|T037|T84.099A|ICD10CM|OTHER MECHANICAL COMPLICATION OF UNSPECIFIED INTERNAL JOINT PROSTHESIS, INITIAL ENCOUNTER|MECH COMPL OF UNSP INTERNAL JOINT PROSTHESIS, INIT ENCNTR
C4083073|T047||ICD10CM|ACUTE SYSTOLIC (CONGESTIVE) HEART FAILURE
C1135191|T047|I50.20|ICD10CM|UNSPECIFIED SYSTOLIC (CONGESTIVE) HEART FAILURE|UNSPECIFIED SYSTOLIC (CONGESTIVE) HEART FAILURE
C2733492|T047||ICD10CM|ACUTE ON CHRONIC SYSTOLIC (CONGESTIVE) HEART FAILURE
C1135194|T047||ICD10CM|CHRONIC SYSTOLIC (CONGESTIVE) HEART FAILURE
C2832062|T037|S06.302A|ICD10CM|UNSPECIFIED FOCAL TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|UNSP FOCAL TBI W LOSS OF CONSCIOUSNESS OF 31-59 MIN, INIT
C2869888|T037|S98.911D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT FOOT, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMP OF RIGHT FOOT, LEVEL UNSP, SUBS
C4269564|T037|S02.672S|ICD10CM|FRACTURE OF ALVEOLUS OF LEFT MANDIBLE, SEQUELA|FRACTURE OF ALVEOLUS OF LEFT MANDIBLE, SEQUELA
C2901198|T046|M84.533A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, RIGHT RADIUS, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, RIGHT RADIUS, INIT
C2869889|T037|S98.911S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT FOOT, LEVEL UNSPECIFIED, SEQUELA|COMPLETE TRAUMATIC AMP OF RIGHT FOOT, LEVEL UNSP, SEQUELA
C4268249|T048|F15.222|ICD10CM|OTHER STIMULANT DEPENDENCE WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE|AMPHETAMINE OR OTHER STIMULANT USE DISORDER, SEVERE, WITH AMPHETAMINE OR OTHER STIMULANT INTOXICATION, WITH PERCEPTUAL DISTURBANCES
C4509229|T047|I50.89|ICD10CM|OTHER HEART FAILURE|OTHER HEART FAILURE
C2874646|T048|F15.220|ICD10CM|OTHER STIMULANT DEPENDENCE WITH INTOXICATION, UNCOMPLICATED|OTHER STIMULANT DEPENDENCE WITH INTOXICATION, UNCOMPLICATED
C2874647|T048|F15.221|ICD10CM|OTHER STIMULANT DEPENDENCE WITH INTOXICATION DELIRIUM|OTHER STIMULANT DEPENDENCE WITH INTOXICATION DELIRIUM
C2895360|T047|M49.89|ICD10CM|SPONDYLOPATHY IN DISEASES CLASSIFIED ELSEWHERE, MULTIPLE SITES IN SPINE|SPOND IN DISEASES CLASSD ELSWHR, MULTIPLE SITES IN SPINE
C4268251|T048|F15.229|ICD10CM|OTHER STIMULANT DEPENDENCE WITH INTOXICATION, UNSPECIFIED|AMPHETAMINE OR OTHER STIMULANT USE DISORDER, SEVERE, WITH AMPHETAMINE OR OTHER STIMULANT INTOXICATION, WITHOUT PERCEPTUAL DISTURBANCES
C2873981|T047|E09.39|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH OTHER DIABETIC OPHTHALMIC COMPLICATION|DRUG/CHEM DIABETES W OTH DIABETIC OPHTHALMIC COMPLICATION
C2853960|T191|C84.40|ICD10CM|PERIPHERAL T-CELL LYMPHOMA, NOT CLASSIFIED, UNSPECIFIED SITE|PERIPHERAL T-CELL LYMPHOMA, NOT CLASSIFIED, UNSPECIFIED SITE
C2873980|T047|E09.36|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH DIABETIC CATARACT|DRUG/CHEM DIABETES MELLITUS W DIABETIC CATARACT
C0409580|T047|M02.9|DMDICD10|REACTIVE ARTHROPATHY, UNSPECIFIED|REAKTIVE ARTHRITIS, NICHT NAEHER BEZEICHNET
C0392097|T033|Z94.4|DMDICD10|LIVER TRANSPLANT STATUS|ZUSTAND NACH LEBERTRANSPLANTATION
C4509307|T047|L97.418|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT HEEL AND MIDFOOT WITH OTHER SPECIFIED SEVERITY|NON-PRS CHRONIC ULCER OF RIGHT HEEL/MIDFT WITH OTH SEVERITY
C0476660|T033|Z94.3|DMDICD10|HEART AND LUNGS TRANSPLANT STATUS|ZUSTAND NACH HERZ-LUNGEN-TRANSPLANTATION
C2889416|T047|M06.219|ICD10CM|RHEUMATOID BURSITIS, UNSPECIFIED SHOULDER|RHEUMATOID BURSITIS, UNSPECIFIED SHOULDER
C0392098|T033|Z94.2|DMDICD10|LUNG TRANSPLANT STATUS|ZUSTAND NACH LUNGENTRANSPLANTATION
C3161075|T047|D61.818|ICD10CM|OTHER PANCYTOPENIA|OTHER PANCYTOPENIA
C0392095|T033|Z94.1|DMDICD10|HEART TRANSPLANT STATUS|ZUSTAND NACH HERZTRANSPLANTATION
C2875346|T047|G83.13|ICD10CM|MONOPLEGIA OF LOWER LIMB AFFECTING RIGHT NONDOMINANT SIDE|MONOPLEGIA OF LOWER LIMB AFFECTING RIGHT NONDOMINANT SIDE
C3161073|T046|D61.810|ICD10CM|ANTINEOPLASTIC CHEMOTHERAPY INDUCED PANCYTOPENIA|ANTINEOPLASTIC CHEMOTHERAPY INDUCED PANCYTOPENIA
C2874639|T048|F15.181|ICD10CM|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED SEXUAL DYSFUNCTION|OTH STIMULANT ABUSE W STIMULANT-INDUCED SEXUAL DYSFUNCTION
C2857342|T037|S72.126A|ICD10CM|NONDISPLACED FRACTURE OF LESSER TROCHANTER OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF LESSER TROCHANTER OF UNSP FEMUR, INIT
C2857343|T037|S72.126B|ICD10CM|NONDISPLACED FRACTURE OF LESSER TROCHANTER OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF LESS TROCHANTER OF UNSP FEMR, 7THB
C2875344|T047|G83.11|ICD10CM|MONOPLEGIA OF LOWER LIMB AFFECTING RIGHT DOMINANT SIDE|MONOPLEGIA OF LOWER LIMB AFFECTING RIGHT DOMINANT SIDE
C2901869|T047|M86.419|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, UNSPECIFIED SHOULDER|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, UNSP SHOULDER
C2874884|T048|F31.32|ICD10CM|BIPOLAR DISORDER, CURRENT EPISODE DEPRESSED, MODERATE|BIPOLAR DISORDER, CURRENT EPISODE DEPRESSED, MODERATE
C0840006|T047|M86.8X8|ICD10CM|OTHER OSTEOMYELITIS, OTHER SITE|OTHER OSTEOMYELITIS, OTHER SITE
C2874882|T048|F31.3|ICD10CM|BIPOLAR DISORDER, CURRENT EPISODE DEPRESSED, MILD OR MODERATE SEVERITY, UNSPECIFIED|BIPOLAR DISORDER, CURRENT EPISODE DEPRESSED, MILD OR MODERATE SEVERITY
C2874883|T048|F31.31|ICD10CM|BIPOLAR DISORDER, CURRENT EPISODE DEPRESSED, MILD|BIPOLAR DISORDER, CURRENT EPISODE DEPRESSED, MILD
C2901867|T047|M86.411|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, RIGHT SHOULDER|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, RIGHT SHOULDER
C2901868|T047|M86.412|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, LEFT SHOULDER|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, LEFT SHOULDER
C0839978|T047|M86.59|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, MULTIPLE SITES|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, MULTIPLE SITES
C2875165|T047|G43.519|ICD10CM|PERSISTENT MIGRAINE AURA WITHOUT CEREBRAL INFARCTION, INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|PERST MIGRAINE AURA W/O CEREBRAL INFRC, NTRCT, W/O STAT MIGR
C2888144|T047|L12.31|ICD10CM|EPIDERMOLYSIS BULLOSA DUE TO DRUG|EPIDERMOLYSIS BULLOSA DUE TO DRUG
C0079293|T047|L12.30|ICD10CM|ACQUIRED EPIDERMOLYSIS BULLOSA, UNSPECIFIED|ACQUIRED EPIDERMOLYSIS BULLOSA, UNSPECIFIED
C2884218|T037|T53.1X2A|ICD10CM|TOXIC EFFECT OF CHLOROFORM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CHLOROFORM, INTENTIONAL SELF-HARM, INIT
C2888145|T047|L12.35|ICD10CM|OTHER ACQUIRED EPIDERMOLYSIS BULLOSA|OTHER ACQUIRED EPIDERMOLYSIS BULLOSA
C2875164|T047|G43.511|ICD10CM|PERSISTENT MIGRAINE AURA WITHOUT CEREBRAL INFARCTION, INTRACTABLE, WITH STATUS MIGRAINOSUS|PERST MIGRAINE AURA W/O CEREBRAL INFRC, NTRCT, W STAT MIGR
C0376358|T191|C61|DMDICD10|MALIGNANT NEOPLASM OF PROSTATE|BOESARTIGE NEUBILDUNG DER PROSTATA
C0840138|T047|M89.60|ICD10AM|OSTEOPATHY AFTER POLIOMYELITIS, UNSPECIFIED SITE|OSTEOPATHY AFTER POLIOMYELITIS, MULTIPLE SITES
C2888784|T047|L98.429|ICD10CM|NON-PRESSURE CHRONIC ULCER OF BACK WITH UNSPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF BACK WITH UNSPECIFIED SEVERITY
C4509343|T047|L98.428|ICD10CM|NON-PRESSURE CHRONIC ULCER OF BACK WITH OTHER SPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF BACK WITH OTH SEVERITY
C2879673|T037|T47.0X2S|ICD10CM|POISONING BY HISTAMINE H2-RECEPTOR BLOCKERS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY HISTAMINE H2-RECEPTOR BLOCKERS, SELF-HARM, SEQUELA
C4509341|T047|L98.425|ICD10CM|NON-PRESSURE CHRONIC ULCER OF BACK WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULCER OF BACK WITH MUSCLE INVL W/O EVD OF NECR
C2888783|T047||ICD10CM|NON-PRESSURE CHRONIC ULCER OF BACK WITH NECROSIS OF BONE
C0078917|T019|E70.319|ICD10CM|OCULAR ALBINISM, UNSPECIFIED|OCULAR ALBINISM, UNSPECIFIED
C2888780|T047|L98.421|ICD10CM|NON-PRESSURE CHRONIC ULCER OF BACK LIMITED TO BREAKDOWN OF SKIN|NON-PRESSURE CHRONIC ULCER OF BACK LIMITED TO BRKDWN SKIN
C2888782|T047||ICD10CM|NON-PRESSURE CHRONIC ULCER OF BACK WITH NECROSIS OF MUSCLE
C2888781|T047||ICD10CM|NON-PRESSURE CHRONIC ULCER OF BACK WITH FAT LAYER EXPOSED
C2889558|T047|M08.232|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, LEFT WRIST|JUVENILE RHEUMATOID ARTHRITIS W SYSTEMIC ONSET, LEFT WRIST
C2889557|T047|M08.231|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, RIGHT WRIST|JUVENILE RHEUMATOID ARTHRITIS W SYSTEMIC ONSET, RIGHT WRIST
C2842025|T191|C46.50|ICD10CM|KAPOSI'S SARCOMA OF UNSPECIFIED LUNG|KAPOSI'S SARCOMA OF UNSPECIFIED LUNG
C2888861|T047|M00.211|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, RIGHT SHOULDER|OTHER STREPTOCOCCAL ARTHRITIS, RIGHT SHOULDER
C2888862|T047|M00.212|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, LEFT SHOULDER|OTHER STREPTOCOCCAL ARTHRITIS, LEFT SHOULDER
C4269272|T037|S02.118A|ICD10CM|OTHER FRACTURE OF OCCIPUT, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTHER FRACTURE OF OCCIPUT, UNSPECIFIED SIDE, INIT
C4269273|T037|S02.118B|ICD10CM|OTHER FRACTURE OF OCCIPUT, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTHER FRACTURE OF OCCIPUT, UNSPECIFIED SIDE, 7THB
C2888863|T047|M00.219|ICD10CM|OTHER STREPTOCOCCAL ARTHRITIS, UNSPECIFIED SHOULDER|OTHER STREPTOCOCCAL ARTHRITIS, UNSPECIFIED SHOULDER
C2835371|T037|S22.060B|ICD10CM|WEDGE COMPRESSION FRACTURE OF T7-T8 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|WEDGE COMPRSN FRACTURE OF T7-T8 VERTEBRA, INIT FOR OPN FX
C2835370|T037|S22.060A|ICD10CM|WEDGE COMPRESSION FRACTURE OF T7-T8 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|WEDGE COMPRESSION FRACTURE OF T7-T8 VERTEBRA, INIT
C2873994|T047|E09.52|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH DIABETIC PERIPHERAL ANGIOPATHY WITH GANGRENE|DRUG/CHEM DIABETES W DIABETIC PRPH ANGIOPATH W GANGRENE
C2905685|T037|X73.2XXS|ICD10CM|INTENTIONAL SELF-HARM BY MACHINE GUN DISCHARGE, SEQUELA|INTENTIONAL SELF-HARM BY MACHINE GUN DISCHARGE, SEQUELA
C2873992|T047|E09.51|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH DIABETIC PERIPHERAL ANGIOPATHY WITHOUT GANGRENE|DRUG/CHEM DIABETES W DIABETIC PRPH ANGIOPATH W/O GANGRENE
C2905683|T037|X73.2XXA|ICD10CM|INTENTIONAL SELF-HARM BY MACHINE GUN DISCHARGE, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY MACHINE GUN DISCHARGE, INIT ENCNTR
C0837024|T047||ICD10CM|TYPE 2 DIABETES MELLITUS WITH KETOACIDOSIS WITH COMA
C0837023|T047||ICD10CM|TYPE 2 DIABETES MELLITUS WITH KETOACIDOSIS WITHOUT COMA
C2855962|T037|S68.421S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT HAND AT WRIST LEVEL, SEQUELA|PARTIAL TRAUMATIC AMP OF RIGHT HAND AT WRIST LEVEL, SEQUELA
C0840001|T047|M86.8X3|ICD10CM|OTHER OSTEOMYELITIS, FOREARM|OTHER OSTEOMYELITIS, FOREARM
C2889209|T047|M05.331|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT WRIST|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF R WRIST
C2876159|T037|T31.74|ICD10CM|BURNS INVOLVING 70-79% OF BODY SURFACE WITH 40-49% THIRD DEGREE BURNS|BURNS OF 70-79% OF BODY SURFACE W 40-49% THIRD DEGREE BURNS
C2876160|T037|T31.75|ICD10CM|BURNS INVOLVING 70-79% OF BODY SURFACE WITH 50-59% THIRD DEGREE BURNS|BURNS OF 70-79% OF BODY SURFACE W 50-59% THIRD DEGREE BURNS
C2876161|T037|T31.76|ICD10CM|BURNS INVOLVING 70-79% OF BODY SURFACE WITH 60-69% THIRD DEGREE BURNS|BURNS OF 70-79% OF BODY SURFACE W 60-69% THIRD DEGREE BURNS
C2876162|T037|T31.77|ICD10CM|BURNS INVOLVING 70-79% OF BODY SURFACE WITH 70-79% THIRD DEGREE BURNS|BURNS OF 70-79% OF BODY SURFACE W 70-79% THIRD DEGREE BURNS
C2837661|T037|S32.10XB|ICD10CM|UNSPECIFIED FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF SACRUM, INIT ENCNTR FOR OPEN FRACTURE
C2855960|T037|S68.421A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT HAND AT WRIST LEVEL, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP OF RIGHT HAND AT WRIST LEVEL, INIT
C2876158|T037|T31.73|ICD10CM|BURNS INVOLVING 70-79% OF BODY SURFACE WITH 30-39% THIRD DEGREE BURNS|BURNS OF 70-79% OF BODY SURFACE W 30-39% THIRD DEGREE BURNS
C2869765|T037|S98.019S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED FOOT AT ANKLE LEVEL, SEQUELA|COMPLETE TRAUMATIC AMP OF UNSP FOOT AT ANKLE LEVEL, SEQUELA
C2883760|T037|T50.902A|ICD10CM|POISONING BY UNSPECIFIED DRUGS, MEDICAMENTS AND BIOLOGICAL SUBSTANCES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY UNSP DRUG/MEDS/BIOL SUBST, SELF-HARM, INIT
C2858338|T037|S72.411A|ICD10CM|DISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED UNSP CONDYLE FX LOWER END OF RIGHT FEMUR, INIT
C2901394|T046|M84.621A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, RIGHT HUMERUS, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, RIGHT HUMERUS, INIT
C2869763|T037|S98.019A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED FOOT AT ANKLE LEVEL, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMP OF UNSP FOOT AT ANKLE LEVEL, INIT
C2858340|T037|S72.411C|ICD10CM|DISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL UNSP CONDYLE FX LOW END R FEMR, 7THC
C2883762|T037|T50.902S|ICD10CM|POISONING BY UNSPECIFIED DRUGS, MEDICAMENTS AND BIOLOGICAL SUBSTANCES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY UNSP DRUG/MEDS/BIOL SUBST, SELF-HARM, SEQUELA
C2883711|T037|T50.7X2S|ICD10CM|POISONING BY ANALEPTICS AND OPIOID RECEPTOR ANTAGONISTS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY ANALEPTICS AND OPIOID RECEPTOR ANTAG, SLF-HRM, SQLA
C2889135|T047|M05.111|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT SHOULDER|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF R SHOULDER
C2895327|T037|M48.54XA|ICD10CM|COLLAPSED VERTEBRA, NOT ELSEWHERE CLASSIFIED, THORACIC REGION, INITIAL ENCOUNTER FOR FRACTURE|COLLAPSED VERTEBRA, NEC, THORACIC REGION, INIT
C2860036|T037|S78.921A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT HIP AND THIGH, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP OF R HIP AND THIGH, LEVEL UNSP, INIT
C2833614|T037|S12.64XB|ICD10CM|TYPE III TRAUMATIC SPONDYLOLISTHESIS OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE III TRAUM SPONDYLOLYSIS OF 7TH CERVCAL VERT, 7THB
C2833613|T037|S12.64XA|ICD10CM|TYPE III TRAUMATIC SPONDYLOLISTHESIS OF SEVENTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE III TRAUM SPONDYLOLYSIS OF SEVENTH CERVCAL VERT, INIT
C2890612|T037|T84.119A|ICD10CM|BREAKDOWN (MECHANICAL) OF INTERNAL FIXATION DEVICE OF UNSPECIFIED BONE OF LIMB, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF INT FIX OF UNSP BONE OF LIMB, INIT
C2890638|T037|T84.125A|ICD10CM|DISPLACEMENT OF INTERNAL FIXATION DEVICE OF LEFT FEMUR, INITIAL ENCOUNTER|DISPLACEMENT OF INTERNAL FIXATION DEVICE OF LEFT FEMUR, INIT
C2890859|T037|T84.620A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL FIXATION DEVICE OF RIGHT FEMUR, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INT FIX OF RIGHT FEMUR, INIT
C2901517|T046|M84.662A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, LEFT TIBIA, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, LEFT TIBIA, INIT
C0839928|T047||ICD10AM|ACUTE HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED SITE
C2832158|T037|S06.325S|ICD10CM|CONTUSION AND LACERATION OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, SEQUELA|CONTUS/LAC L CEREB W LOC >24 HR W RET CONSC LEV, SEQUELA
C2860037|T037|S78.921D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT HIP AND THIGH, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMP OF R HIP AND THIGH, LEVEL UNSP, SUBS
C0839936|T047||ICD10AM|ACUTE HEMATOGENOUS OSTEOMYELITIS, OTHER SITES
C0839928|T047|M86.09|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, MULTIPLE SITES|ACUTE HEMATOGENOUS OSTEOMYELITIS, MULTIPLE SITES
C0263369|T047|L94.5|DMDICD10|RETIFORM PARAPSORIASIS|POIKILODERMIA ATROPHICANS VASCULARIS [JACOBI]
C0162442|T047|L41.4|DMDICD10|LARGE PLAQUE PARAPSORIASIS|GROSSFLECKIGE PARAPSORIASIS EN PLAQUES
C0263370|T047|L41.3|DMDICD10|SMALL PLAQUE PARAPSORIASIS|KLEINFLECKIGE PARAPSORIASIS EN PLAQUES
C0162851|T047|L41.1|DMDICD10|PITYRIASIS LICHENOIDES CHRONICA|PARAPSORIASIS GUTTATA
C0162852|T047|L41.0|DMDICD10|PITYRIASIS LICHENOIDES ET VARIOLIFORMIS ACUTA|PITYRIASIS LICHENOIDES ET VARIOLIFORMIS ACUTA [MUCHA-HABERMANN]
C2832156|T037|S06.325A|ICD10CM|CONTUSION AND LACERATION OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, INITIAL ENCOUNTER|CONTUS/LAC LEFT CEREBRUM W LOC >24 HR W RET CONSC LEV, INIT
C0030491|T047|L41.9|DMDICD10|PARAPSORIASIS, UNSPECIFIED|PARAPSORIASIS, NICHT NAEHER BEZEICHNET
C0477486|T047|L41.8|DMDICD10|OTHER PARAPSORIASIS|SONSTIGE PARAPSORIASIS
C0477324|T047|D81.89|ICD10CM|OTHER COMBINED IMMUNODEFICIENCIES|OTHER COMBINED IMMUNODEFICIENCIES
C2882415|T047|I63.59|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF OTHER CEREBRAL ARTERY|CEREB INFRC DUE TO UNSP OCCLS OR STENOSIS OF CEREBRAL ARTERY
C2887822|T047|K51.50|ICD10CM|LEFT SIDED COLITIS WITHOUT COMPLICATIONS|LEFT SIDED COLITIS WITHOUT COMPLICATIONS
C2858644|T037|S72.441A|ICD10CM|DISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF LOWER EPIPHYSIS (SEPARATION) OF RIGHT FEMUR, INIT
C2891134|T037|T85.611D|ICD10CM|BREAKDOWN (MECHANICAL) OF INTRAPERITONEAL DIALYSIS CATHETER, SUBSEQUENT ENCOUNTER|BREAKDOWN OF INTRAPERITONEAL DIALYSIS CATHETER, SUBS
C2891133|T037|T85.611A|ICD10CM|BREAKDOWN (MECHANICAL) OF INTRAPERITONEAL DIALYSIS CATHETER, INITIAL ENCOUNTER|BREAKDOWN OF INTRAPERITONEAL DIALYSIS CATHETER, INIT
C0155970|T047|K25.1|DMDICD10|ACUTE GASTRIC ULCER WITH PERFORATION|ULCUS VENTRICULI: AKUT, MIT PERFORATION
C0155973|T047|K25.2|DMDICD10|ACUTE GASTRIC ULCER WITH BOTH HEMORRHAGE AND PERFORATION|ULCUS VENTRICULI: AKUT, MIT BLUTUNG UND PERFORATION
C0155982|T047|K25.5|DMDICD10|CHRONIC OR UNSPECIFIED GASTRIC ULCER WITH PERFORATION|ULCUS VENTRICULI: CHRONISCH ODER NICHT NAEHER BEZEICHNET, MIT PERFORATION
C2889093|T047|M02.849|ICD10CM|OTHER REACTIVE ARTHROPATHIES, UNSPECIFIED HAND|OTHER REACTIVE ARTHROPATHIES, UNSPECIFIED HAND
C2889092|T047|M02.842|ICD10CM|OTHER REACTIVE ARTHROPATHIES, LEFT HAND|OTHER REACTIVE ARTHROPATHIES, LEFT HAND
C2889091|T047|M02.841|ICD10CM|OTHER REACTIVE ARTHROPATHIES, RIGHT HAND|OTHER REACTIVE ARTHROPATHIES, RIGHT HAND
C2882402|T047|I63.519|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF UNSPECIFIED MIDDLE CEREBRAL ARTERY|CEREB INFRC D/T UNSP OCCLS OR STENOS OF UNSP MID CEREB ART
C2856760|T037|S72.035C|ICD10CM|NONDISPLACED MIDCERVICAL FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP MIDCERVICAL FX L FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2882400|T047|I63.511|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF RIGHT MIDDLE CEREBRAL ARTERY|CEREB INFRC D/T UNSP OCCLS OR STENOS OF RIGHT MID CEREB ART
C2882401|T047|I63.512|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF LEFT MIDDLE CEREBRAL ARTERY|CEREB INFRC D/T UNSP OCCLS OR STENOS OF LEFT MID CEREB ART
C4268489|T047|I63.513|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF BILATERAL MIDDLE CEREBRAL ARTERIES|CEREB INFRC D/T UNSP OCCLS OR STENOS OF BI MIDDLE CEREB ART
C2833301|T037|S12.190A|ICD10CM|OTHER DISPLACED FRACTURE OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH DISP FX OF SECOND CERVICAL VERTEBRA, INIT FOR CLOS FX
C2833510|T037|S12.491B|ICD10CM|OTHER NONDISPLACED FRACTURE OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH NONDISP FX OF FIFTH CERVICAL VERTEBRA, INIT FOR OPN FX
C2833509|T037|S12.491A|ICD10CM|OTHER NONDISPLACED FRACTURE OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH NONDISP FX OF FIFTH CERVICAL VERTEBRA, INIT FOR CLOS FX
C2890410|T037|T84.012A|ICD10CM|BROKEN INTERNAL RIGHT KNEE PROSTHESIS, INITIAL ENCOUNTER|BROKEN INTERNAL RIGHT KNEE PROSTHESIS, INITIAL ENCOUNTER
C2890550|T037|T84.069A|ICD10CM|WEAR OF ARTICULAR BEARING SURFACE OF UNSPECIFIED INTERNAL PROSTHETIC JOINT, INITIAL ENCOUNTER|WEAR OF ARTIC BEARING SURFACE OF UNSP INT PROSTH JOINT, INIT
C0155995|T047|K26.1|DMDICD10|ACUTE DUODENAL ULCER WITH PERFORATION|ULCUS DUODENI: AKUT, MIT PERFORATION
C0868862|T047|M46.1|DMDICD10|SACROILIITIS, NOT ELSEWHERE CLASSIFIED|SAKROILIITIS, ANDERENORTS NICHT KLASSIFIZIERT
C0840047|T046|M87.38|ICD10AM|OTHER SECONDARY OSTEONECROSIS, OTHER SITE|OTHER SECONDARY OSTEONECROSIS, OTHER SITE
C0342751|T047||ICD10CM|POMPE DISEASE
C2837553|T037|S32.030A|ICD10CM|WEDGE COMPRESSION FRACTURE OF THIRD LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|WEDGE COMPRESSION FRACTURE OF THIRD LUMBAR VERTEBRA, INIT
C2837554|T037|S32.030B|ICD10CM|WEDGE COMPRESSION FRACTURE OF THIRD LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|WEDGE COMPRSN FX THIRD LUM VERTEBRA, INIT FOR OPN FX
C4267995|T047|E09.3543|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, BILATERAL|DRUG/CHEM DIAB WITH PROLIF DIAB RTNOP WITH COMB DETACH, BI
C4267994|T047|E09.3542|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, LEFT EYE|DRUG/CHEM DIAB W PROLIF DIAB RTNOP WITH COMB DETACH, L EYE
C4267993|T047|E09.3541|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, RIGHT EYE|DRUG/CHEM DIAB W PROLIF DIAB RTNOP WITH COMB DETACH, R EYE
C2837525|T037|S32.021B|ICD10CM|STABLE BURST FRACTURE OF SECOND LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|STABLE BURST FX SECOND LUM VERTEBRA, INIT FOR OPN FX
C2837524|T037|S32.021A|ICD10CM|STABLE BURST FRACTURE OF SECOND LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|STABLE BURST FRACTURE OF SECOND LUMBAR VERTEBRA, INIT
C4267996|T047|E09.3549|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, UNSPECIFIED EYE|DRUG/CHEM DIAB WITH PROLIF DIAB RTNOP WITH COMB DETACH, UNSP
C2886724|T037|T79.1XXA|ICD10CM|FAT EMBOLISM (TRAUMATIC), INITIAL ENCOUNTER|FAT EMBOLISM (TRAUMATIC), INITIAL ENCOUNTER
C2876621|T037|T36.3X2S|ICD10CM|POISONING BY MACROLIDES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY MACROLIDES, INTENTIONAL SELF-HARM, SEQUELA
C2882634|T047|I69.861|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING RIGHT DOMINANT SIDE|OTH PARLYT SYND FOL OTH CEREBVASC DISEASE AFF RIGHT DOM SIDE
C2902126|T046|M87.81|ICD10CM|OTHER OSTEONECROSIS, UNSPECIFIED SHOULDER|OTHER OSTEONECROSIS, SHOULDER
C2858712|T037|S72.445A|ICD10CM|NONDISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF LOWER EPIPHYSIS (SEPARATION) OF L FEMUR, INIT
C2858713|T037|S72.445B|ICD10CM|NONDISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF LOW EPIPHY (SEPARATION) OF L FEMR, 7THB
C2858714|T037|S72.445C|ICD10CM|NONDISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF LOW EPIPHY (SEPARATION) OF L FEMR, 7THC
C2902128|T046|M87.812|ICD10CM|OTHER OSTEONECROSIS, LEFT SHOULDER|OTHER OSTEONECROSIS, LEFT SHOULDER
C2902127|T046|M87.811|ICD10CM|OTHER OSTEONECROSIS, RIGHT SHOULDER|OTHER OSTEONECROSIS, RIGHT SHOULDER
C2837795|T037|S32.2XXA|ICD10CM|FRACTURE OF COCCYX, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF COCCYX, INITIAL ENCOUNTER FOR CLOSED FRACTURE
C2837796|T037|S32.2XXB|ICD10CM|FRACTURE OF COCCYX, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF COCCYX, INITIAL ENCOUNTER FOR OPEN FRACTURE
C4270491|T046|T85.123A|ICD10CM|DISPLACEMENT OF IMPLANTED ELECTRONIC NEUROSTIMULATOR, GENERATOR, INITIAL ENCOUNTER|DISPLACEMENT OF IMPLNT ELEC NSTIM, GENERATOR, INIT
C2856003|T037|S68.610S|ICD10CM|COMPLETE TRAUMATIC TRANSPHALANGEAL AMPUTATION OF RIGHT INDEX FINGER, SEQUELA|COMPLETE TRAUMATIC TRNSPHAL AMP OF R IDX FNGR, SEQUELA
C2882175|T047|I25.701|ICD10CM|ATHEROSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT(S), UNSPECIFIED, WITH ANGINA PECTORIS WITH DOCUMENTED SPASM|ATHSCL CABG, UNSP, W ANGINA PECTORIS W DOCUMENTED SPASM
C2882174|T047|I25.700|ICD10CM|ATHEROSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT(S), UNSPECIFIED, WITH UNSTABLE ANGINA PECTORIS|ATHEROSCLEROSIS OF CABG, UNSP, W UNSTABLE ANGINA PECTORIS
C2838000|T191|C43.70|ICD10CM|MALIGNANT MELANOMA OF UNSPECIFIED LOWER LIMB, INCLUDING HIP|MALIGNANT MELANOMA OF UNSPECIFIED LOWER LIMB, INCLUDING HIP
C2838001|T191|C43.71|ICD10CM|MALIGNANT MELANOMA OF RIGHT LOWER LIMB, INCLUDING HIP|MALIGNANT MELANOMA OF RIGHT LOWER LIMB, INCLUDING HIP
C2838002|T191|C43.72|ICD10CM|MALIGNANT MELANOMA OF LEFT LOWER LIMB, INCLUDING HIP|MALIGNANT MELANOMA OF LEFT LOWER LIMB, INCLUDING HIP
C2882177|T047|I25.709|ICD10CM|ATHEROSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT(S), UNSPECIFIED, WITH UNSPECIFIED ANGINA PECTORIS|ATHEROSCLEROSIS OF CABG, UNSP, W UNSP ANGINA PECTORIS
C2882176|T047|I25.708|ICD10CM|ATHEROSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT(S), UNSPECIFIED, WITH OTHER FORMS OF ANGINA PECTORIS|ATHEROSCLEROSIS OF CABG, UNSP, W OTH ANGINA PECTORIS
C2885852|T037|T63.792S|ICD10CM|TOXIC EFFECT OF CONTACT WITH OTHER VENOMOUS PLANT, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CONTACT W OTH VENOM PLANT, SLF-HRM, SEQUELA
C2854041|T191|C85.28|ICD10CM|MEDIASTINAL (THYMIC) LARGE B-CELL LYMPHOMA, LYMPH NODES OF MULTIPLE SITES|MEDIASTINAL (THYMIC) LARGE B-CELL LYMPHOMA, NODES MULT SITE
C2886210|T037|T65.92XS|ICD10CM|TOXIC EFFECT OF UNSPECIFIED SUBSTANCE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF UNSP SUBSTANCE, SELF-HARM, SEQUELA
C2889926|T037|T82.328A|ICD10CM|DISPLACEMENT OF OTHER VASCULAR GRAFTS, INITIAL ENCOUNTER|DISPLACEMENT OF OTHER VASCULAR GRAFTS, INITIAL ENCOUNTER
C2885850|T037|T63.792A|ICD10CM|TOXIC EFFECT OF CONTACT WITH OTHER VENOMOUS PLANT, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CONTACT W OTH VENOMOUS PLANT, SLF-HRM, INIT
C2848391|T037|S58.011S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT ELBOW LEVEL, RIGHT ARM, SEQUELA|COMPLETE TRAUMATIC AMP AT ELBOW LEVEL, RIGHT ARM, SEQUELA
C2859993|T037|S78.029D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT UNSPECIFIED HIP JOINT, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION AT UNSP HIP JOINT, SUBS ENCNTR
C0153809|T191||ICD10CM|MYCOSIS FUNGOIDES, LYMPH NODES OF MULTIPLE SITES
C2853956|T191|C84.09|ICD10CM|MYCOSIS FUNGOIDES, EXTRANODAL AND SOLID ORGAN SITES|MYCOSIS FUNGOIDES, EXTRANODAL AND SOLID ORGAN SITES
C2848389|T037|S58.011A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT ELBOW LEVEL, RIGHT ARM, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMP AT ELBOW LEVEL, RIGHT ARM, INIT
C0153803|T191||ICD10CM|MYCOSIS FUNGOIDES, INTRATHORACIC LYMPH NODES
C0153804|T191||ICD10CM|MYCOSIS FUNGOIDES, INTRA-ABDOMINAL LYMPH NODES
C0026948|T191|C84.00|ICD10CM|MYCOSIS FUNGOIDES, UNSPECIFIED SITE|MYCOSIS FUNGOIDES, UNSPECIFIED SITE
C0153802|T191|C84.01|ICD10CM|MYCOSIS FUNGOIDES, LYMPH NODES OF HEAD, FACE, AND NECK|MYCOSIS FUNGOIDES, LYMPH NODES OF HEAD, FACE, AND NECK
C0153807|T191||ICD10CM|MYCOSIS FUNGOIDES, INTRAPELVIC LYMPH NODES
C0153808|T191||ICD10CM|MYCOSIS FUNGOIDES, SPLEEN
C0153805|T191|C84.04|ICD10CM|MYCOSIS FUNGOIDES, LYMPH NODES OF AXILLA AND UPPER LIMB|MYCOSIS FUNGOIDES, LYMPH NODES OF AXILLA AND UPPER LIMB
C0153806|T191|C84.05|ICD10CM|MYCOSIS FUNGOIDES, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|MYCOSIS FUNGOIDES, NODES OF INGUINAL REGION AND LOWER LIMB
C2888801|T047|M00.029|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, UNSPECIFIED ELBOW|STAPHYLOCOCCAL ARTHRITIS, UNSPECIFIED ELBOW
C2835284|T037|S22.038B|ICD10CM|OTHER FRACTURE OF THIRD THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF THIRD THORACIC VERTEBRA, INIT FOR OPN FX
C2835283|T037|S22.038A|ICD10CM|OTHER FRACTURE OF THIRD THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF THIRD THORACIC VERTEBRA, INIT FOR CLOS FX
C2888800|T047|M00.022|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, LEFT ELBOW|STAPHYLOCOCCAL ARTHRITIS, LEFT ELBOW
C2888799|T047|M00.021|ICD10CM|STAPHYLOCOCCAL ARTHRITIS, RIGHT ELBOW|STAPHYLOCOCCAL ARTHRITIS, RIGHT ELBOW
C2859992|T037|S78.029A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT UNSPECIFIED HIP JOINT, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION AT UNSP HIP JOINT, INIT ENCNTR
C2882834|T047|I70.442|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF CALF|ATHSCL AUTOL VEIN BYPASS OF THE LEFT LEG W ULCER OF CALF
C2882835|T047|I70.443|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF ANKLE|ATHSCL AUTOL VEIN BYPASS OF THE LEFT LEG W ULCER OF ANKLE
C2882833|T047|I70.441|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF THIGH|ATHSCL AUTOL VEIN BYPASS OF THE LEFT LEG W ULCER OF THIGH
C2882837|T047|I70.444|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF HEEL AND MIDFOOT|ATHSCL AUTOL VEIN BYPASS OF LEFT LEG W ULC OF HEEL AND MIDFT
C2882839|T047|I70.445|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF OTHER PART OF FOOT|ATHSCL AUTOL VEIN BYPASS OF LEFT LEG W ULCER OTH PRT FOOT
C4269315|T037|S02.11FB|ICD10CM|TYPE III OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE III OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, 7THB
C2882840|T047|I70.448|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF OTHER PART OF LOWER LEG|ATHSCL AUTOL VEIN BYPASS OF LEFT LEG W ULCER OTH PRT LOW LEG
C3648033|T191|C82.65|ICD10CM|CUTANEOUS FOLLICLE CENTER LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|CUTAN FOLICL CNTR LYMPH, NODES OF ING REGION AND LOWER LIMB
C2832026|T037|S06.2X3S|ICD10CM|DIFFUSE TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, SEQUELA|DIFFUSE TBI W LOC OF 1-5 HRS 59 MIN, SEQUELA
C4269314|T037|S02.11FA|ICD10CM|TYPE III OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE III OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, INIT
C2832024|T037|S06.2X3A|ICD10CM|DIFFUSE TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|DIFFUSE TBI W LOSS OF CONSCIOUSNESS OF 1-5 HRS 59 MIN, INIT
C2832008|T037|S06.1X9A|ICD10CM|TRAUMATIC CEREBRAL EDEMA WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|TRAUMATIC CEREBRAL EDEMA W LOC OF UNSP DURATION, INIT
C2874709|T048|F16.920|ICD10CM|HALLUCINOGEN USE, UNSPECIFIED WITH INTOXICATION, UNCOMPLICATED|HALLUCINOGEN USE, UNSP WITH INTOXICATION, UNCOMPLICATED
C2883359|T037|T49.3X2S|ICD10CM|POISONING BY EMOLLIENTS, DEMULCENTS AND PROTECTANTS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY EMOLLIENTS, DEMULCENTS AND PROTECT, SLF-HRM, SQLA
C2832010|T037|S06.1X9S|ICD10CM|TRAUMATIC CEREBRAL EDEMA WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|TRAUMATIC CEREBRAL EDEMA W LOC OF UNSP DURATION, SEQUELA
C2874515|T048|F13.12|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE WITH INTOXICATION, UNSPECIFIED|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE WITH INTOXICATION
C2855846|T037|S68.019S|ICD10CM|COMPLETE TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF UNSPECIFIED THUMB, SEQUELA|COMPLETE TRAUMATIC MCP AMPUTATION OF THMB, SEQUELA
C2883357|T037|T49.3X2A|ICD10CM|POISONING BY EMOLLIENTS, DEMULCENTS AND PROTECTANTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY EMOLLIENTS, DEMULCENTS AND PROTECT, SELF-HARM, INIT
C2874514|T048|F13.121|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE WITH INTOXICATION DELIRIUM|SEDATV/HYP/ANXIOLYTC ABUSE W INTOXICATION DELIRIUM
C2874519|T048|F13.151|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC ABUSE WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|SEDATV/HYP/ANXIOLYTC ABUSE W PSYCHOTIC DISORDER W HALLUCIN
C2842121|T191|C50.619|ICD10CM|MALIGNANT NEOPLASM OF AXILLARY TAIL OF UNSPECIFIED FEMALE BREAST|MALIGNANT NEOPLASM OF AXILLARY TAIL OF UNSP FEMALE BREAST
C2842120|T191|C50.612|ICD10CM|MALIGNANT NEOPLASM OF AXILLARY TAIL OF LEFT FEMALE BREAST|MALIGNANT NEOPLASM OF AXILLARY TAIL OF LEFT FEMALE BREAST
C2842119|T191|C50.611|ICD10CM|MALIGNANT NEOPLASM OF AXILLARY TAIL OF RIGHT FEMALE BREAST|MALIGNANT NEOPLASM OF AXILLARY TAIL OF RIGHT FEMALE BREAST
C2833887|T037|S14.112D|ICD10CM|COMPLETE LESION AT C2 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION AT C2 LEVEL OF CERVICAL SPINAL CORD, SUBS
C2833886|T037|S14.112A|ICD10CM|COMPLETE LESION AT C2 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION AT C2 LEVEL OF CERVICAL SPINAL CORD, INIT
C2861578|T191||ICD10CM|ACUTE MYELOBLASTIC LEUKEMIA, IN RELAPSE
C0153886|T191||ICD10CM|ACUTE MYELOBLASTIC LEUKEMIA, IN REMISSION
C2861577|T191||ICD10CM|ACUTE MYELOBLASTIC LEUKEMIA, NOT HAVING ACHIEVED REMISSION
C2833888|T037|S14.112S|ICD10CM|COMPLETE LESION AT C2 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|COMPLETE LESION AT C2 LEVEL OF CERVICAL SPINAL CORD, SEQUELA
C2865570|T037|S88.911S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT LOWER LEG, LEVEL UNSPECIFIED, SEQUELA|COMPLETE TRAUMATIC AMP OF R LOW LEG, LEVEL UNSP, SEQUELA
C4269319|T037|S02.11FS|ICD10CM|TYPE III OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, SEQUELA|TYPE III OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, SEQUELA
C2877973|T037|T41.3X2S|ICD10CM|POISONING BY LOCAL ANESTHETICS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY LOCAL ANESTHETICS, SELF-HARM, SEQUELA
C2889412|T047|M06.08|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, VERTEBRAE|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, VERTEBRAE
C2889413|T047|M06.09|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, MULTIPLE SITES|RHEUMATOID ARTHRITIS W/O RHEUMATOID FACTOR, MULTIPLE SITES
C2832276|T037|S06.353S|ICD10CM|TRAUMATIC HEMORRHAGE OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 1 HOURS TO 5 HOURS 59 MINUTES, SEQUELA|TRAUM HEMOR L CEREB W LOC OF 1-5 HRS 59 MINUTES, SEQUELA
C2889387|T047|M06.00|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, UNSPECIFIED SITE|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, UNSP SITE
C2877971|T037|T41.3X2A|ICD10CM|POISONING BY LOCAL ANESTHETICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY LOCAL ANESTHETICS, INTENTIONAL SELF-HARM, INIT
C2832395|T037|S06.382A|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF BRAINSTEM WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|CONTUS/LAC/HEM BRAINSTEM W LOC OF 31-59 MIN, INIT
C2832274|T037|S06.353A|ICD10CM|TRAUMATIC HEMORRHAGE OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 1 HOURS TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|TRAUM HEMOR LEFT CEREBRUM W LOC OF 1-5 HRS 59 MINUTES, INIT
C2886756|T037|T79.A12A|ICD10CM|TRAUMATIC COMPARTMENT SYNDROME OF LEFT UPPER EXTREMITY, INITIAL ENCOUNTER|TRAUMATIC COMPARTMENT SYNDROME OF LEFT UPPER EXTREMITY, INIT
C2889628|T047|M08.912|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, LEFT SHOULDER|JUVENILE ARTHRITIS, UNSPECIFIED, LEFT SHOULDER
C2889627|T047|M08.911|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, RIGHT SHOULDER|JUVENILE ARTHRITIS, UNSPECIFIED, RIGHT SHOULDER
C2889629|T047|M08.919|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, UNSPECIFIED SHOULDER|JUVENILE ARTHRITIS, UNSPECIFIED, UNSPECIFIED SHOULDER
C2837890|T037|S32.401A|ICD10CM|UNSPECIFIED FRACTURE OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF RIGHT ACETABULUM, INIT FOR CLOS FX
C2837891|T037|S32.401B|ICD10CM|UNSPECIFIED FRACTURE OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF RIGHT ACETABULUM, INIT FOR OPN FX
C4268114|T047|E11.3553|ICD10CM|TYPE 2 DIABETES MELLITUS WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, BILATERAL|TYPE 2 DIABETES WITH STABLE PROLIF DIABETIC RTNOP, BILATERAL
C4268113|T047|E11.3552|ICD10CM|TYPE 2 DIABETES MELLITUS WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, LEFT EYE|TYPE 2 DIABETES WITH STABLE PROLIF DIABETIC RTNOP, LEFT EYE
C4268112|T047|E11.3551|ICD10CM|TYPE 2 DIABETES MELLITUS WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, RIGHT EYE|TYPE 2 DIABETES WITH STABLE PROLIF DIABETIC RTNOP, RIGHT EYE
C0393949|T047|I67.89|ICD10CM|OTHER CEREBROVASCULAR DISEASE|OTHER CEREBROVASCULAR DISEASE
C0026708|T047||ICD10CM|SCHEIE'S SYNDROME
C0086431|T047||ICD10CM|HURLER-SCHEIE SYNDROME
C4268115|T047|E11.3559|ICD10CM|TYPE 2 DIABETES MELLITUS WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, UNSPECIFIED EYE|TYPE 2 DIABETES WITH STABLE PROLIF DIABETIC RTNOP, UNSP
C3264376|T047|I67.81|ICD10CM|ACUTE CEREBROVASCULAR INSUFFICIENCY|ACUTE CEREBROVASCULAR INSUFFICIENCY UNSPECIFIED AS TO LOCATION OR REVERSIBILITY
C0917798|T047||ICD10CM|CEREBRAL ISCHEMIA
C2910843|T033|Z44.112|ICD10CM|ENCOUNTER FOR FITTING AND ADJUSTMENT OF COMPLETE LEFT ARTIFICIAL LEG|ENCOUNTER FOR FIT/ADJST OF COMPLETE LEFT ARTIFICIAL LEG
C2910842|T033|Z44.111|ICD10CM|ENCOUNTER FOR FITTING AND ADJUSTMENT OF COMPLETE RIGHT ARTIFICIAL LEG|ENCOUNTER FOR FIT/ADJST OF COMPLETE RIGHT ARTIFICIAL LEG
C2910844|T033|Z44.119|ICD10CM|ENCOUNTER FOR FITTING AND ADJUSTMENT OF COMPLETE ARTIFICIAL LEG, UNSPECIFIED LEG|ENCOUNTER FOR FIT/ADJST OF COMPLETE ARTIFICIAL LEG, UNSP LEG
C2874482|T048|F12.19|ICD10CM|CANNABIS ABUSE WITH UNSPECIFIED CANNABIS-INDUCED DISORDER|CANNABIS ABUSE WITH UNSPECIFIED CANNABIS-INDUCED DISORDER
C0477416|T047|G90.8|DMDICD10|OTHER DISORDERS OF AUTONOMIC NERVOUS SYSTEM|SONSTIGE KRANKHEITEN DES AUTONOMEN NERVENSYSTEMS
C1145628|T047|G90|DMDICD10|DISORDER OF THE AUTONOMIC NERVOUS SYSTEM, UNSPECIFIED|KRANKHEITEN DES AUTONOMEN NERVENSYSTEMS
C2835774|T037|S24.109S|ICD10CM|UNSPECIFIED INJURY AT UNSPECIFIED LEVEL OF THORACIC SPINAL CORD, SEQUELA|UNSP INJURY AT UNSP LEVEL OF THORACIC SPINAL CORD, SEQUELA
C2890019|T037|T82.515A|ICD10CM|BREAKDOWN (MECHANICAL) OF UMBRELLA DEVICE, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF UMBRELLA DEVICE, INITIAL ENCOUNTER
C3264370|T046|I48.3|ICD10CM|TYPICAL ATRIAL FLUTTER|TYPICAL ATRIAL FLUTTER
C0013364|T047|G90.1|DMDICD10|FAMILIAL DYSAUTONOMIA [RILEY-DAY]|FAMILIAERE DYSAUTONOMIE [RILEY-DAY-SYNDROM]
C0865487|T047|G90.2|ICD10CM|HORNER'S SYNDROME|CERVICAL SYMPATHETIC DYSTROPHY OR PARALYSIS
C0235480|T047|I48.0|ICD10CM|PAROXYSMAL ATRIAL FIBRILLATION|PAROXYSMAL ATRIAL FIBRILLATION
C0238015|T047||ICD10CM|AUTONOMIC DYSREFLEXIA
C3264372|T033|I48.4|ICD10CM|ATYPICAL ATRIAL FLUTTER|ATYPICAL ATRIAL FLUTTER
C2874011|T047|E09.649|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH HYPOGLYCEMIA WITHOUT COMA|DRUG/CHEM DIABETES MELLITUS W HYPOGLYCEMIA W/O COMA
C2874010|T047|E09.641|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH HYPOGLYCEMIA WITH COMA|DRUG/CHEM DIABETES MELLITUS W HYPOGLYCEMIA W COMA
C2911415|T033|Z89.432|ICD10CM|ACQUIRED ABSENCE OF LEFT FOOT|ACQUIRED ABSENCE OF LEFT FOOT
C2884625|T037|T56.92XA|ICD10CM|TOXIC EFFECT OF UNSPECIFIED METAL, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF UNSP METAL, INTENTIONAL SELF-HARM, INIT
C2910346|T047|Q87.418|ICD10CM|MARFAN'S SYNDROME WITH OTHER CARDIOVASCULAR MANIFESTATIONS|MARFAN'S SYNDROME WITH OTHER CARDIOVASCULAR MANIFESTATIONS
C2886119|T037|T65.6X2A|ICD10CM|TOXIC EFFECT OF PAINTS AND DYES, NOT ELSEWHERE CLASSIFIED, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF PAINTS AND DYES, NEC, SELF-HARM, INIT
C2910345|T047|Q87.410|ICD10CM|MARFAN'S SYNDROME WITH AORTIC DILATION|MARFAN'S SYNDROME WITH AORTIC DILATION
C0040021|T047|I73.1|DMDICD10|THROMBOANGIITIS OBLITERANS [BUERGER'S DISEASE]|THROMBANGIITIS OBLITERANS [ENDANGIITIS VON-WINIWARTER-BUERGER]
C2911414|T033|Z89.431|ICD10CM|ACQUIRED ABSENCE OF RIGHT FOOT|ACQUIRED ABSENCE OF RIGHT FOOT
C2884627|T037|T56.92XS|ICD10CM|TOXIC EFFECT OF UNSPECIFIED METAL, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF UNSP METAL, INTENTIONAL SELF-HARM, SEQUELA
C0085617|T046|I73.9|ICD10CM|PERIPHERAL VASCULAR DISEASE, UNSPECIFIED|SPASM OF ARTERY
C2886121|T037|T65.6X2S|ICD10CM|TOXIC EFFECT OF PAINTS AND DYES, NOT ELSEWHERE CLASSIFIED, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF PAINTS AND DYES, NEC, SELF-HARM, SEQUELA
C0155763|T047|I77.8|ICD10CM|OTHER SPECIFIED DISORDERS OF ARTERIES AND ARTERIOLES|OTHER SPECIFIED DISORDERS OF ARTERIES AND ARTERIOLES
C2884723|T037|T57.92XS|ICD10CM|TOXIC EFFECT OF UNSPECIFIED INORGANIC SUBSTANCE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF UNSP INORGANIC SUBSTANCE, SELF-HARM, SEQUELA
C0037773|T047|G11.4|DMDICD10|HEREDITARY SPASTIC PARAPLEGIA|HEREDITAERE SPASTISCHE PARAPLEGIE
C2874191|T047|E24.0|ICD10CM|PITUITARY-DEPENDENT CUSHING'S DISEASE|OVERPRODUCTION OF PITUITARY ACTH
C4268956|T046|N99.532|ICD10CM|MALFUNCTION OF CONTINENT STOMA OF URINARY TRACT|MALFUNCTION OF CONTINENT STOMA OF URINARY TRACT
C4268957|T046|N99.533|ICD10CM|HERNIATION OF CONTINENT STOMA OF URINARY TRACT|HERNIATION OF CONTINENT STOMA OF URINARY TRACT
C4268954|T046|N99.530|ICD10CM|HEMORRHAGE OF CONTINENT STOMA OF URINARY TRACT|HEMORRHAGE OF CONTINENT STOMA OF URINARY TRACT
C4268955|T046|N99.531|ICD10CM|INFECTION OF CONTINENT STOMA OF URINARY TRACT|INFECTION OF CONTINENT STOMA OF URINARY TRACT
C4268958|T046|N99.534|ICD10CM|STENOSIS OF CONTINENT STOMA OF URINARY TRACT|STENOSIS OF CONTINENT STOMA OF URINARY TRACT
C0481241|T037|Y62.2|DMDICD10|FAILURE OF STERILE PRECAUTIONS DURING KIDNEY DIALYSIS AND OTHER PERFUSION|UNZULAENGLICHE ASEPTISCHE KAUTELEN: BEI HAEMODIALYSE ODER SONSTIGER PERFUSION
C4268959|T046|N99.538|ICD10CM|OTHER COMPLICATION OF CONTINENT STOMA OF URINARY TRACT|OTHER COMPLICATION OF CONTINENT STOMA OF URINARY TRACT
C0024776|T047|E71.0|DMDICD10|MAPLE-SYRUP-URINE DISEASE|AHORNSIRUP- (HARN-) KRANKHEIT
C2911416|T033|Z89.439|ICD10CM|ACQUIRED ABSENCE OF UNSPECIFIED FOOT|ACQUIRED ABSENCE OF UNSPECIFIED FOOT
C2889145|T047|M05.132|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT WRIST|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889144|T047|M05.131|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT WRIST|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF R WRIST
C2889146|T047|M05.139|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP WRIST
C2882695|T047|I70.208|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES, OTHER EXTREMITY|UNSP ATHSCL NATIVE ARTERIES OF EXTREMITIES, OTH EXTREMITY
C2882696|T047|I70.209|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES, UNSPECIFIED EXTREMITY|UNSP ATHSCL NATIVE ARTERIES OF EXTREMITIES, UNSP EXTREMITY
C2977876|T037|S32.599A|ICD10CM|OTHER SPECIFIED FRACTURE OF UNSPECIFIED PUBIS, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF UNSP PUBIS, INIT ENCNTR FOR CLOSED FRACTURE
C2910224|T047||ICD10CM|CYSTIC DILATATION OF COLLECTING DUCTS
C2874066|T047|E10.630|ICD10CM|TYPE 1 DIABETES MELLITUS WITH PERIODONTAL DISEASE|TYPE 1 DIABETES MELLITUS WITH PERIODONTAL DISEASE
C2882692|T047|I70.201|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES, RIGHT LEG|UNSP ATHSCL NATIVE ARTERIES OF EXTREMITIES, RIGHT LEG
C2882693|T047|I70.202|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES, LEFT LEG|UNSP ATHSCL NATIVE ARTERIES OF EXTREMITIES, LEFT LEG
C2882694|T047|I70.203|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES, BILATERAL LEGS|UNSP ATHSCL NATIVE ARTERIES OF EXTREMITIES, BILATERAL LEGS
C2910225|T047|Q61.19|ICD10CM|OTHER POLYCYSTIC KIDNEY, INFANTILE TYPE|OTHER POLYCYSTIC KIDNEY, INFANTILE TYPE
C2874067|T047|E10.638|ICD10CM|TYPE 1 DIABETES MELLITUS WITH OTHER ORAL COMPLICATIONS|TYPE 1 DIABETES MELLITUS WITH OTHER ORAL COMPLICATIONS
C2887779|T047|K50.90|ICD10CM|CROHN'S DISEASE, UNSPECIFIED, WITHOUT COMPLICATIONS|CROHN'S DISEASE, UNSPECIFIED, WITHOUT COMPLICATIONS
C4268612|T047|K55.012|ICD10CM|DIFFUSE ACUTE (REVERSIBLE) ISCHEMIA OF SMALL INTESTINE|DIFFUSE ACUTE (REVERSIBLE) ISCHEMIA OF SMALL INTESTINE
C2874446|T048|F11.251|ICD10CM|OPIOID DEPENDENCE WITH OPIOID-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|OPIOID DEPEND W OPIOID-INDUC PSYCHOTIC DISORDER W HALLUCIN
C2874445|T048|F11.250|ICD10CM|OPIOID DEPENDENCE WITH OPIOID-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|OPIOID DEPEND W OPIOID-INDUC PSYCHOTIC DISORDER W DELUSIONS
C2890132|T037|T82.7XXA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO OTHER CARDIAC AND VASCULAR DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|INFECT/INFLM REACT D/T OTH CARDI/VASC DEV/IMPLNT/GRFT, INIT
C2858217|T037|S72.366B|ICD10CM|NONDISPLACED SEGMENTAL FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP SEG FX SHAFT OF UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2858218|T037|S72.366C|ICD10CM|NONDISPLACED SEGMENTAL FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP SEG FX SHAFT OF UNSP FEMR, 7THC
C2874447|T048|F11.259|ICD10CM|OPIOID DEPENDENCE WITH OPIOID-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|OPIOID DEPENDENCE WITH OPIOID-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED
C4268613|T047|K55.019|ICD10CM|ACUTE (REVERSIBLE) ISCHEMIA OF SMALL INTESTINE, EXTENT UNSPECIFIED|ACUTE ISCHEMIA OF SMALL INTESTINE, EXTENT UNSPECIFIED
C2876720|T037|T36.7X2S|ICD10CM|POISONING BY ANTIFUNGAL ANTIBIOTICS, SYSTEMICALLY USED, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ANTIFUNG ANTIBIOT, SYS USED, SELF-HARM, SEQUELA
C2856569|T037|S72.019B|ICD10CM|UNSPECIFIED INTRACAPSULAR FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP INTRACAP FX UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2869829|T037|S98.149D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF ONE UNSPECIFIED LESSER TOE, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF ONE UNSP LESSER TOE, SUBS
C2835162|T037|S22.001B|ICD10CM|STABLE BURST FRACTURE OF UNSPECIFIED THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|STABLE BURST FRACTURE OF UNSP THOR VERTEBRA, INIT FOR OPN FX
C2835161|T037|S22.001A|ICD10CM|STABLE BURST FRACTURE OF UNSPECIFIED THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|STABLE BURST FRACTURE OF UNSP THORACIC VERTEBRA, INIT
C2874761|T048|F18.221|ICD10CM|INHALANT DEPENDENCE WITH INTOXICATION DELIRIUM|INHALANT DEPENDENCE WITH INTOXICATION DELIRIUM
C0153379|T191|C06.2|DMDICD10|MALIGNANT NEOPLASM OF RETROMOLAR AREA|BOESARTIGE NEUBILDUNG: RETROMOLARREGION
C2833839|T191|C06.1|ICD10CM|MALIGNANT NEOPLASM OF VESTIBULE OF MOUTH|MALIGNANT NEOPLASM OF LABIAL SULCUS (UPPER) (LOWER)
C2833837|T191|C06.0|ICD10CM|MALIGNANT NEOPLASM OF CHEEK MUCOSA|MALIGNANT NEOPLASM OF INTERNAL CHEEK
C0864852|T191|C06.9|ICD10CM|MALIGNANT NEOPLASM OF MOUTH, UNSPECIFIED|MALIGNANT NEOPLASM OF MINOR SALIVARY GLAND, UNSPECIFIED SITE
C2902082|T046|M87.311|ICD10CM|OTHER SECONDARY OSTEONECROSIS, RIGHT SHOULDER|OTHER SECONDARY OSTEONECROSIS, RIGHT SHOULDER
C2902083|T046|M87.312|ICD10CM|OTHER SECONDARY OSTEONECROSIS, LEFT SHOULDER|OTHER SECONDARY OSTEONECROSIS, LEFT SHOULDER
C2900968|T046|M84.444A|ICD10CM|PATHOLOGICAL FRACTURE, RIGHT FINGER(S), INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, RIGHT FINGER(S), INIT FOR FX
C2900925|T046|M84.433A|ICD10CM|PATHOLOGICAL FRACTURE, RIGHT RADIUS, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, RIGHT RADIUS, INIT FOR FX
C4270181|T046|T82.868A|ICD10CM|THROMBOSIS DUE TO VASCULAR PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|THROMBOSIS DUE TO VASCULAR PROSTH DEV/GRFT, INIT
C2869901|T037|S98.921D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT FOOT, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF RIGHT FOOT, LEVEL UNSP, SUBS
C2837495|T037|S32.012A|ICD10CM|UNSTABLE BURST FRACTURE OF FIRST LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSTABLE BURST FRACTURE OF FIRST LUMBAR VERTEBRA, INIT
C2905744|T037|X77.8XXS|ICD10CM|INTENTIONAL SELF-HARM BY OTHER HOT OBJECTS, SEQUELA|INTENTIONAL SELF-HARM BY OTHER HOT OBJECTS, SEQUELA
C2837496|T037|S32.012B|ICD10CM|UNSTABLE BURST FRACTURE OF FIRST LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSTABLE BURST FX FIRST LUM VERTEBRA, INIT FOR OPN FX
C4270451|T046|T85.110A|ICD10CM|BREAKDOWN (MECHANICAL) OF IMPLANTED ELECTRONIC NEUROSTIMULATOR OF BRAIN ELECTRODE (LEAD), INITIAL ENCOUNTER|BREAKDOWN OF IMPLNT ELEC NSTIM OF BRAIN LEAD, INIT
C1299613|T047|E10.8|DMDICD10|TYPE 1 DIABETES MELLITUS WITH UNSPECIFIED COMPLICATIONS|PRIMAER INSULINABHAENGIGER DIABETES MELLITUS [TYP-I-DIABETES]: MIT NICHT NAEHER BEZEICHNETEN KOMPLIKATIONEN
C0494284|T047|E10.9|DMDICD10|TYPE 1 DIABETES MELLITUS WITHOUT COMPLICATIONS|PRIMAER INSULINABHAENGIGER DIABETES MELLITUS [TYP-I-DIABETES]: OHNE KOMPLIKATIONEN
C4269531|T037|S02.651A|ICD10CM|FRACTURE OF ANGLE OF RIGHT MANDIBLE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF ANGLE OF RIGHT MANDIBLE, INIT
C2838207|T037|S32.455A|ICD10CM|NONDISPLACED TRANSVERSE FRACTURE OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED TRANSVERSE FRACTURE OF LEFT ACETABULUM, INIT
C2888614|T047|L89.899|ICD10CM|PRESSURE ULCER OF OTHER SITE, UNSPECIFIED STAGE|PRESSURE ULCER OF OTHER SITE, UNSPECIFIED STAGE
C2900526|T046|M80.861A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, RIGHT LOWER LEG, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, R LOW LEG, INIT
C2888605|T047|L89.892|ICD10CM|PRESSURE ULCER OF OTHER SITE, STAGE 2|PRESSURE ULCER OF OTHER SITE, STAGE 2
C2888608|T047|L89.893|ICD10CM|PRESSURE ULCER OF OTHER SITE, STAGE 3|PRESSURE ULCER OF OTHER SITE, STAGE 3
C2888599|T047|L89.890|ICD10CM|PRESSURE ULCER OF OTHER SITE, UNSTAGEABLE|PRESSURE ULCER OF OTHER SITE, UNSTAGEABLE
C2888602|T047|L89.891|ICD10CM|PRESSURE ULCER OF OTHER SITE, STAGE 1|PRESSURE ULCER OF OTHER SITE, STAGE 1
C4269277|T037|S02.118S|ICD10CM|OTHER FRACTURE OF OCCIPUT, UNSPECIFIED SIDE, SEQUELA|OTHER FRACTURE OF OCCIPUT, UNSPECIFIED SIDE, SEQUELA
C2888611|T047|L89.894|ICD10CM|PRESSURE ULCER OF OTHER SITE, STAGE 4|PRESSURE ULCER OF OTHER SITE, STAGE 4
C2857615|T037|S72.24XA|ICD10CM|NONDISPLACED SUBTROCHANTERIC FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED SUBTROCHANTERIC FRACTURE OF RIGHT FEMUR, INIT
C2857617|T037|S72.24XC|ICD10CM|NONDISPLACED SUBTROCHANTERIC FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP SUBTROCHNT FX R FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2857616|T037|S72.24XB|ICD10CM|NONDISPLACED SUBTROCHANTERIC FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP SUBTROCHNT FX RIGHT FEMUR, INIT FOR OPN FX TYPE I/2
C2905800|T037|X82.2XXS|ICD10CM|INTENTIONAL COLLISION OF MOTOR VEHICLE WITH TREE, SEQUELA|INTENTIONAL COLLISION OF MOTOR VEHICLE WITH TREE, SEQUELA
C2832710|T037|S06.9X9S|ICD10CM|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|UNSP INTRACRANIAL INJURY W LOC OF UNSP DURATION, SEQUELA
C2835442|T037|S22.080A|ICD10CM|WEDGE COMPRESSION FRACTURE OF T11-T12 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|WEDGE COMPRESSION FRACTURE OF T11-T12 VERTEBRA, INIT
C2874456|T048|F11.921|ICD10CM|OPIOID USE, UNSPECIFIED WITH INTOXICATION DELIRIUM|OPIOID USE, UNSPECIFIED WITH INTOXICATION DELIRIUM
C2874455|T048|F11.920|ICD10CM|OPIOID USE, UNSPECIFIED WITH INTOXICATION, UNCOMPLICATED|OPIOID USE, UNSPECIFIED WITH INTOXICATION, UNCOMPLICATED
C2874457|T048|F11.922|ICD10CM|OPIOID USE, UNSPECIFIED WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE|OPIOID USE, UNSP W INTOXICATION WITH PERCEPTUAL DISTURBANCE
C2838394|T037|S32.519B|ICD10CM|FRACTURE OF SUPERIOR RIM OF UNSPECIFIED PUBIS, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF SUPERIOR RIM OF UNSP PUBIS, INIT FOR OPN FX
C2905798|T037|X82.2XXA|ICD10CM|INTENTIONAL COLLISION OF MOTOR VEHICLE WITH TREE, INITIAL ENCOUNTER|INTENTIONAL COLLISION OF MOTOR VEHICLE W TREE, INIT ENCNTR
C2832708|T037|S06.9X9A|ICD10CM|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|UNSP INTRACRANIAL INJURY W LOC OF UNSP DURATION, INIT
C2874458|T048|F11.929|ICD10CM|OPIOID USE, UNSPECIFIED WITH INTOXICATION, UNSPECIFIED|OPIOID USE, UNSPECIFIED WITH INTOXICATION, UNSPECIFIED
C2833205|T037|S12.091B|ICD10CM|OTHER NONDISPLACED FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH NONDISP FX OF FIRST CERVICAL VERTEBRA, INIT FOR OPN FX
C2833204|T037|S12.091A|ICD10CM|OTHER NONDISPLACED FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH NONDISP FX OF FIRST CERVICAL VERTEBRA, INIT FOR CLOS FX
C2905799|T037|X82.2XXD|ICD10CM|INTENTIONAL COLLISION OF MOTOR VEHICLE WITH TREE, SUBSEQUENT ENCOUNTER|INTENTIONAL COLLISION OF MOTOR VEHICLE W TREE, SUBS ENCNTR
C2887196|T047|I83.028|ICD10CM|VARICOSE VEINS OF LEFT LOWER EXTREMITY WITH ULCER OTHER PART OF LOWER LEG|VARICOSE VEINS OF L LOW EXTREM W ULCER OTH PART OF LOWER LEG
C2887197|T047|I83.029|ICD10CM|VARICOSE VEINS OF LEFT LOWER EXTREMITY WITH ULCER OF UNSPECIFIED SITE|VARICOSE VEINS OF LEFT LOWER EXTREMITY W ULCER OF UNSP SITE
C2861636|T191||ICD10CM|MAST CELL LEUKEMIA NOT HAVING ACHIEVED REMISSION
C0836977|T191||ICD10AM|MAST CELL LEUKEMIA, IN REMISSION
C2367254|T191||ICD10CM|MAST CELL LEUKEMIA, IN RELAPSE
C2887195|T047|I83.025|ICD10CM|VARICOSE VEINS OF LEFT LOWER EXTREMITY WITH ULCER OTHER PART OF FOOT|VARICOSE VEINS OF L LOW EXTREM W ULCER OTH PART OF FOOT
C2887190|T047|I83.022|ICD10CM|VARICOSE VEINS OF LEFT LOWER EXTREMITY WITH ULCER OF CALF|VARICOSE VEINS OF LEFT LOWER EXTREMITY WITH ULCER OF CALF
C2887191|T047|I83.023|ICD10CM|VARICOSE VEINS OF LEFT LOWER EXTREMITY WITH ULCER OF ANKLE|VARICOSE VEINS OF LEFT LOWER EXTREMITY WITH ULCER OF ANKLE
C2860200|T037|S79.139A|ICD10CM|SALTER-HARRIS TYPE III PHYSEAL FRACTURE OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SLTR-HARIS TYPE III PHYSEAL FX LOWER END OF UNSP FEMUR, INIT
C2887189|T047|I83.021|ICD10CM|VARICOSE VEINS OF LEFT LOWER EXTREMITY WITH ULCER OF THIGH|VARICOSE VEINS OF LEFT LOWER EXTREMITY WITH ULCER OF THIGH
C2893633|T047|M12.021|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], RIGHT ELBOW|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], RIGHT ELBOW
C2893634|T047|M12.022|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], LEFT ELBOW|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], LEFT ELBOW
C4270656|T046|T85.890A|ICD10CM|OTHER SPECIFIED COMPLICATION OF NERVOUS SYSTEM PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|OTH COMPLICATION OF NERVOUS SYSTEM PROSTH DEV/GRFT, INIT
C2869799|T037|S98.122D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT GREAT TOE, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF LEFT GREAT TOE, SUBS ENCNTR
C2893635|T047|M12.029|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], UNSPECIFIED ELBOW|CHRONIC POSTRHEUMATIC ARTHROPATHY, UNSPECIFIED ELBOW
C2869798|T037|S98.122A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT GREAT TOE, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF LEFT GREAT TOE, INIT ENCNTR
C2885409|T037|T63.072S|ICD10CM|TOXIC EFFECT OF VENOM OF OTHER AUSTRALIAN SNAKE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF AUSTRALIAN SNAKE, SLF-HRM, SEQUELA
C2837582|T037|S32.039B|ICD10CM|UNSPECIFIED FRACTURE OF THIRD LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF THIRD LUMBAR VERTEBRA, INIT FOR OPN FX
C2869800|T037|S98.122S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT GREAT TOE, SEQUELA|PARTIAL TRAUMATIC AMPUTATION OF LEFT GREAT TOE, SEQUELA
C2874874|T048|F31.10|ICD10CM|BIPOLAR DISORDER, CURRENT EPISODE MANIC WITHOUT PSYCHOTIC FEATURES, UNSPECIFIED|BIPOLAR DISORDER, CURRENT EPISODE MANIC WITHOUT PSYCHOTIC FEATURES, UNSPECIFIED
C2874875|T048|F31.11|ICD10CM|BIPOLAR DISORDER, CURRENT EPISODE MANIC WITHOUT PSYCHOTIC FEATURES, MILD|BIPOLAR DISORD, CRNT EPISODE MANIC W/O PSYCH FEATURES, MILD
C2874876|T048|F31.12|ICD10CM|BIPOLAR DISORDER, CURRENT EPISODE MANIC WITHOUT PSYCHOTIC FEATURES, MODERATE|BIPOLAR DISORD, CRNT EPISODE MANIC W/O PSYCH FEATURES, MOD
C2874877|T048|F31.13|ICD10CM|BIPOLAR DISORDER, CURRENT EPISODE MANIC WITHOUT PSYCHOTIC FEATURES, SEVERE|BIPOLAR DISORD, CRNT EPSD MANIC W/O PSYCH FEATURES, SEVERE
C2877512|T037|T39.8X2A|ICD10CM|POISONING BY OTHER NONOPIOID ANALGESICS AND ANTIPYRETICS, NOT ELSEWHERE CLASSIFIED, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY OTH NONOPIO ANALGES/ANTIPYRET, NEC, SELF-HARM, INIT
C2882467|T047|I69.054|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING LEFT NON-DOMINANT SIDE|HEMIPLGA FOLLOWING NTRM SUBARACH HEMOR AFF LEFT NONDOM SIDE
C2882466|T047|I69.053|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING RIGHT NON-DOMINANT SIDE|HEMIPLGA FOLLOWING NTRM SUBARACH HEMOR AFF RIGHT NONDOM SIDE
C2882465|T047|I69.052|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING LEFT DOMINANT SIDE|HEMIPLGA FOL NTRM SUBARACH HEMOR AFF LEFT DOMINANT SIDE
C2882464|T047|I69.051|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING RIGHT DOMINANT SIDE|HEMIPLGA FOL NTRM SUBARACH HEMOR AFF RIGHT DOMINANT SIDE
C2837876|T037|S32.392B|ICD10CM|OTHER FRACTURE OF LEFT ILIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTHER FRACTURE OF LEFT ILIUM, INIT ENCNTR FOR OPEN FRACTURE
C2857309|T037|S72.124B|ICD10CM|NONDISPLACED FRACTURE OF LESSER TROCHANTER OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF LESS TROCHANTER OF R FEMR, 7THB
C2857310|T037|S72.124C|ICD10CM|NONDISPLACED FRACTURE OF LESSER TROCHANTER OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF LESS TROCHANTER OF R FEMR, 7THC
C2857308|T037|S72.124A|ICD10CM|NONDISPLACED FRACTURE OF LESSER TROCHANTER OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF LESSER TROCHANTER OF RIGHT FEMUR, INIT
C2882468|T047|I69.059|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING UNSPECIFIED SIDE|HEMIPLGA FOLLOWING NTRM SUBARACH HEMOR AFFECTING UNSP SIDE
C2886474|T037|T71.232A|ICD10CM|ASPHYXIATION DUE TO BEING TRAPPED IN A (DISCARDED) REFRIGERATOR, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|ASPHYX D/T BEING TRAP IN A (DISCARDED) REFRIG, SLF-HRM, INIT
C2905675|T037|X73.0XXA|ICD10CM|INTENTIONAL SELF-HARM BY SHOTGUN DISCHARGE, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY SHOTGUN DISCHARGE, INIT ENCNTR
C2838266|T037|S32.471B|ICD10CM|DISPLACED FRACTURE OF MEDIAL WALL OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISP FX OF MEDIAL WALL OF RIGHT ACETABULUM, INIT FOR OPN FX
C2838265|T037|S32.471A|ICD10CM|DISPLACED FRACTURE OF MEDIAL WALL OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF MEDIAL WALL OF RIGHT ACETABULUM, INIT FOR CLOS FX
C2905676|T037|X73.0XXD|ICD10CM|INTENTIONAL SELF-HARM BY SHOTGUN DISCHARGE, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY SHOTGUN DISCHARGE, SUBS ENCNTR
C2886476|T037|T71.232S|ICD10CM|ASPHYXIATION DUE TO BEING TRAPPED IN A (DISCARDED) REFRIGERATOR, INTENTIONAL SELF-HARM, SEQUELA|ASPHYX D/T BEING TRAP IN A (DISCARDED) REFRIG, SLF-HRM, SQLA
C2882163|T047|I25.110|ICD10CM|ATHEROSCLEROTIC HEART DISEASE OF NATIVE CORONARY ARTERY WITH UNSTABLE ANGINA PECTORIS|ATHSCL HEART DISEASE OF NATIVE COR ART W UNSTABLE ANG PCTRS
C2882164|T047|I25.111|ICD10CM|ATHEROSCLEROTIC HEART DISEASE OF NATIVE CORONARY ARTERY WITH ANGINA PECTORIS WITH DOCUMENTED SPASM|ATHSCL HEART DISEASE OF NATIVE COR ART W ANG PCTRS W SPASM
C2837446|T037|S32.000B|ICD10CM|WEDGE COMPRESSION FRACTURE OF UNSPECIFIED LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|WEDGE COMPRSN FRACTURE OF UNSP LUM VERTEBRA, INIT FOR OPN FX
C2837445|T037|S32.000A|ICD10CM|WEDGE COMPRESSION FRACTURE OF UNSPECIFIED LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|WEDGE COMPRESSION FRACTURE OF UNSP LUMBAR VERTEBRA, INIT
C2882165|T047|I25.118|ICD10CM|ATHEROSCLEROTIC HEART DISEASE OF NATIVE CORONARY ARTERY WITH OTHER FORMS OF ANGINA PECTORIS|ATHSCL HEART DISEASE OF NATIVE COR ART W OTH ANG PCTRS
C2882168|T047|I25.119|ICD10CM|ATHEROSCLEROTIC HEART DISEASE OF NATIVE CORONARY ARTERY WITH UNSPECIFIED ANGINA PECTORIS|ATHSCL HEART DISEASE OF NATIVE COR ART W UNSP ANG PCTRS
C2911428|T033|Z89.619|ICD10CM|ACQUIRED ABSENCE OF UNSPECIFIED LEG ABOVE KNEE|ACQUIRED ABSENCE OF UNSPECIFIED LEG ABOVE KNEE
C4269354|T037|S02.32XS|ICD10CM|FRACTURE OF ORBITAL FLOOR, LEFT SIDE, SEQUELA|FRACTURE OF ORBITAL FLOOR, LEFT SIDE, SEQUELA
C4270647|T046|T85.860A|ICD10CM|THROMBOSIS DUE TO NERVOUS SYSTEM PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|THROMBOSIS DUE TO NERVOUS SYSTEM PROSTH DEV/GRFT, INIT
C2830469|T047|R65.20|ICD10CM|SEVERE SEPSIS WITHOUT SEPTIC SHOCK|SEVERE SEPSIS WITHOUT SEPTIC SHOCK
C2830470|T047|R65.21|ICD10CM|SEVERE SEPSIS WITH SEPTIC SHOCK|SEVERE SEPSIS WITH SEPTIC SHOCK
C2883071|T047|I80.229|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF UNSPECIFIED POPLITEAL VEIN|PHLEBITIS AND THROMBOPHLEBITIS OF UNSPECIFIED POPLITEAL VEIN
C4269350|T037|S02.32XB|ICD10CM|FRACTURE OF ORBITAL FLOOR, LEFT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF ORBITAL FLOOR, LEFT SIDE, 7THB
C0265080|T047|I62.00|ICD10CM|NONTRAUMATIC SUBDURAL HEMORRHAGE, UNSPECIFIED|NONTRAUMATIC SUBDURAL HEMORRHAGE, UNSPECIFIED
C0494607|T046||ICD10CM|NONTRAUMATIC ACUTE SUBDURAL HEMORRHAGE
C2882326|T047|I62.02|ICD10CM|NONTRAUMATIC SUBACUTE SUBDURAL HEMORRHAGE|NONTRAUMATIC SUBACUTE SUBDURAL HEMORRHAGE
C2882327|T047|I62.03|ICD10CM|NONTRAUMATIC CHRONIC SUBDURAL HEMORRHAGE|NONTRAUMATIC CHRONIC SUBDURAL HEMORRHAGE
C2883068|T047|I80.221|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF RIGHT POPLITEAL VEIN|PHLEBITIS AND THROMBOPHLEBITIS OF RIGHT POPLITEAL VEIN
C2883070|T047|I80.223|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF POPLITEAL VEIN, BILATERAL|PHLEBITIS AND THROMBOPHLEBITIS OF POPLITEAL VEIN, BILATERAL
C2883069|T047|I80.222|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF LEFT POPLITEAL VEIN|PHLEBITIS AND THROMBOPHLEBITIS OF LEFT POPLITEAL VEIN
C4270463|T046|T85.112A|ICD10CM|BREAKDOWN (MECHANICAL) OF IMPLANTED ELECTRONIC NEUROSTIMULATOR OF SPINAL CORD ELECTRODE (LEAD), INITIAL ENCOUNTER|BREAKDOWN OF IMPLNT ELEC NSTIM OF SPINAL CORD LEAD, INIT
C2889553|T047|M08.21|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, UNSPECIFIED SHOULDER|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, SHOULDER
C4269553|T037|S02.671B|ICD10CM|FRACTURE OF ALVEOLUS OF RIGHT MANDIBLE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF ALVEOLUS OF RIGHT MANDIBLE, 7THB
C2889551|T047|M08.211|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, RIGHT SHOULDER|JUVENILE RHEUMATOID ARTHRITIS W SYSTEMIC ONSET, R SHOULDER
C2889552|T047|M08.212|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, LEFT SHOULDER|JUVENILE RHEUMATOID ARTHRITIS W SYSTEMIC ONSET, L SHOULDER
C4269557|T037|S02.671S|ICD10CM|FRACTURE OF ALVEOLUS OF RIGHT MANDIBLE, SEQUELA|FRACTURE OF ALVEOLUS OF RIGHT MANDIBLE, SEQUELA
C2833190|T037|S12.041B|ICD10CM|NONDISPLACED LATERAL MASS FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP LATERAL MASS FX FIRST CERVCAL VERT, INIT FOR OPN FX
C2832612|T037|S06.825S|ICD10CM|INJURY OF LEFT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, SEQUELA|INJ L INT CRTD, INTCR W LOC >24 HR W RET CONSC LEV, SEQUELA
C2856534|T037|S72.011A|ICD10CM|UNSPECIFIED INTRACAPSULAR FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP INTRACAPSULAR FRACTURE OF RIGHT FEMUR, INIT FOR CLOS FX
C2856536|T037|S72.011C|ICD10CM|UNSPECIFIED INTRACAPSULAR FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP INTRACAP FX RIGHT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2856535|T037|S72.011B|ICD10CM|UNSPECIFIED INTRACAPSULAR FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP INTRACAP FX RIGHT FEMUR, INIT FOR OPN FX TYPE I/2
C2856516|T037|S72.009A|ICD10CM|FRACTURE OF UNSPECIFIED PART OF NECK OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF UNSP PART OF NECK OF UNSP FEMUR, INIT
C2857016|T037|S72.065A|ICD10CM|NONDISPLACED ARTICULAR FRACTURE OF HEAD OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED ARTICULAR FRACTURE OF HEAD OF LEFT FEMUR, INIT
C0837040|T047|E11.36|ICD10AM|TYPE 2 DIABETES MELLITUS WITH DIABETIC CATARACT|TYPE 2 DIABETES MELLITUS WITH DIABETIC CATARACT
C2874096|T047|E11.39|ICD10CM|TYPE 2 DIABETES MELLITUS WITH OTHER DIABETIC OPHTHALMIC COMPLICATION|TYPE 2 DIABETES W OTH DIABETIC OPHTHALMIC COMPLICATION
C2856517|T037|S72.009B|ICD10CM|FRACTURE OF UNSPECIFIED PART OF NECK OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|FX UNSP PART OF NECK OF UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2901778|T047|M86.032|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, LEFT RADIUS AND ULNA|ACUTE HEMATOGENOUS OSTEOMYELITIS, LEFT RADIUS AND ULNA
C2901777|T047|M86.031|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, RIGHT RADIUS AND ULNA|ACUTE HEMATOGENOUS OSTEOMYELITIS, RIGHT RADIUS AND ULNA
C2876129|T037|T31.11|ICD10CM|BURNS INVOLVING 10-19% OF BODY SURFACE WITH 10-19% THIRD DEGREE BURNS|BURNS OF 10-19% OF BODY SURFACE W 10-19% THIRD DEGREE BURNS
C2901779|T047|M86.039|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED RADIUS AND ULNA|ACUTE HEMATOGENOUS OSTEOMYELITIS, UNSP RADIUS AND ULNA
C0496938|T191|D43.4|DMDICD10|NEOPLASM OF UNCERTAIN BEHAVIOR OF SPINAL CORD|NEUBILDUNG UNSICHEREN ODER UNBEKANNTEN VERHALTENS: RUECKENMARK
C2873703|T191||ICD10CM|NEOPLASM OF UNCERTAIN BEHAVIOR OF BRAIN, INFRATENTORIAL
C2873701|T191||ICD10CM|NEOPLASM OF UNCERTAIN BEHAVIOR OF BRAIN, SUPRATENTORIAL
C0496937|T191|D43.3|DMDICD10|NEOPLASM OF UNCERTAIN BEHAVIOR OF CRANIAL NERVES|NEUBILDUNG UNSICHEREN ODER UNBEKANNTEN VERHALTENS: HIRNNERVEN
C2873704|T191|D43.2|ICD10CM|NEOPLASM OF UNCERTAIN BEHAVIOR OF BRAIN, UNSPECIFIED|NEOPLASM OF UNCERTAIN BEHAVIOR OF BRAIN, UNSPECIFIED
C2886394|T037|T71.152A|ICD10CM|ASPHYXIATION DUE TO SMOTHERING IN FURNITURE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|ASPHYXIATION DUE TO SMOTHERING IN FURNITURE, SELF-HARM, INIT
C2873706|T191|D43.9|ICD10CM|NEOPLASM OF UNCERTAIN BEHAVIOR OF CENTRAL NERVOUS SYSTEM, UNSPECIFIED|NEOPLASM OF UNCERTAIN BEHAVIOR OF CNSL, UNSP
C2976850|T191|D43.8|ICD10CM|NEOPLASM OF UNCERTAIN BEHAVIOR OF OTHER SPECIFIED PARTS OF CENTRAL NERVOUS SYSTEM|NEOPLASM OF UNCERTAIN BEHAVIOR OF PRT CENTRAL NERVOUS SYSTEM
C2865555|T037|S88.121A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, RIGHT LOWER LEG, INITIAL ENCOUNTER|PART TRAUM AMP AT LEVEL BETW KNEE AND ANKLE, R LOW LEG, INIT
C2865556|T037|S88.121D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, RIGHT LOWER LEG, SUBSEQUENT ENCOUNTER|PART TRAUM AMP AT LEVEL BETW KNEE AND ANKLE, R LOW LEG, SUBS
C2890064|T037|T82.530A|ICD10CM|LEAKAGE OF SURGICALLY CREATED ARTERIOVENOUS FISTULA, INITIAL ENCOUNTER|LEAKAGE OF SURGICALLY CREATED ARTERIOVENOUS FISTULA, INIT
C2911427|T033|Z89.612|ICD10CM|ACQUIRED ABSENCE OF LEFT LEG ABOVE KNEE|ACQUIRED ABSENCE OF LEFT LEG ABOVE KNEE
C0477617|T047|M48.8|ICD10CM|OTHER SPECIFIED SPONDYLOPATHIES, SITE UNSPECIFIED|OTHER SPECIFIED SPONDYLOPATHIES
C0838677|T047|M48.8X8|ICD10CM|OTHER SPECIFIED SPONDYLOPATHIES, SACRAL AND SACROCOCCYGEAL REGION|OTH SPONDYLOPATHIES, SACRAL AND SACROCOCCYGEAL REGION
C2860016|T037|S78.122S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN LEFT HIP AND KNEE, SEQUELA|PARTIAL TRAUM AMP AT LEVEL BETW LEFT HIP AND KNEE, SEQUELA
C0838674|T047|M48.8X5|ICD10CM|OTHER SPECIFIED SPONDYLOPATHIES, THORACOLUMBAR REGION|OTHER SPECIFIED SPONDYLOPATHIES, THORACOLUMBAR REGION
C0838673|T047|M48.8X4|ICD10CM|OTHER SPECIFIED SPONDYLOPATHIES, THORACIC REGION|OTHER SPECIFIED SPONDYLOPATHIES, THORACIC REGION
C0838676|T047|M48.8X7|ICD10CM|OTHER SPECIFIED SPONDYLOPATHIES, LUMBOSACRAL REGION|OTHER SPECIFIED SPONDYLOPATHIES, LUMBOSACRAL REGION
C0838675|T047|M48.8X6|ICD10CM|OTHER SPECIFIED SPONDYLOPATHIES, LUMBAR REGION|OTHER SPECIFIED SPONDYLOPATHIES, LUMBAR REGION
C0838670|T047|M48.8X1|ICD10CM|OTHER SPECIFIED SPONDYLOPATHIES, OCCIPITO-ATLANTO-AXIAL REGION|OTH SPONDYLOPATHIES, OCCIPITO-ATLANTO-AXIAL REGION
C0838672|T047|M48.8X3|ICD10CM|OTHER SPECIFIED SPONDYLOPATHIES, CERVICOTHORACIC REGION|OTHER SPECIFIED SPONDYLOPATHIES, CERVICOTHORACIC REGION
C0838671|T047|M48.8X2|ICD10CM|OTHER SPECIFIED SPONDYLOPATHIES, CERVICAL REGION|OTHER SPECIFIED SPONDYLOPATHIES, CERVICAL REGION
C2888698|T047|L97.402|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED HEEL AND MIDFOOT WITH FAT LAYER EXPOSED|NON-PRS CHR ULCER OF UNSP HEEL AND MIDFOOT W FAT LAYER EXPOS
C2888699|T047|L97.403|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED HEEL AND MIDFOOT WITH NECROSIS OF MUSCLE|NON-PRS CHR ULCER OF UNSP HEEL AND MIDFOOT W NECROS MUSCLE
C2888697|T047|L97.401|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED HEEL AND MIDFOOT LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHR ULCER OF UNSP HEEL AND MIDFT LMT TO BRKDWN SKIN
C4509303|T047|L97.406|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED HEEL AND MIDFOOT WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC UNSP HEEL/MIDFT W BNE INVL W/O EVD OF NECR
C2888700|T047|L97.404|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED HEEL AND MIDFOOT WITH NECROSIS OF BONE|NON-PRS CHRONIC ULCER OF UNSP HEEL AND MIDFOOT W NECROS BONE
C4509302|T047|L97.405|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED HEEL AND MIDFOOT WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC UNSP HEEL/MIDFT W MSL INVL W/O EVD OF NECR
C2890867|T037|T84.622A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL FIXATION DEVICE OF RIGHT TIBIA, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INT FIX OF RIGHT TIBIA, INIT
C4509304|T047|L97.408|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED HEEL AND MIDFOOT WITH OTHER SPECIFIED SEVERITY|NON-PRS CHRONIC ULCER OF UNSP HEEL/MIDFT WITH OTH SEVERITY
C2888701|T047|L97.409|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED HEEL AND MIDFOOT WITH UNSPECIFIED SEVERITY|NON-PRS CHRONIC ULCER OF UNSP HEEL AND MIDFOOT W UNSP SEVERT
C2977002|T047|I82.502|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF LEFT LOWER EXTREMITY|CHRONIC EMBOLISM AND THOMBOS UNSP DEEP VEINS OF L LOW EXTREM
C2977003|T047|I82.503|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF LOWER EXTREMITY, BILATERAL|CHRONIC EMBLSM AND THOMBOS UNSP DEEP VEINS OF LOW EXTRM, BI
C2901991|T046|M87.12|ICD10CM|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED HUMERUS|OSTEONECROSIS DUE TO DRUGS, HUMERUS
C2977001|T047|I82.501|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF RIGHT LOWER EXTREMITY|CHRONIC EMBOLISM AND THOMBOS UNSP DEEP VEINS OF R LOW EXTREM
C0839956|T047|M86.28|ICD10AM|SUBACUTE OSTEOMYELITIS, OTHER SITE|SUBACUTE OSTEOMYELITIS, OTHER SITE
C0839948|T047|M86.29|ICD10CM|SUBACUTE OSTEOMYELITIS, MULTIPLE SITES|SUBACUTE OSTEOMYELITIS, MULTIPLE SITES
C2901990|T046|M87.122|ICD10CM|OSTEONECROSIS DUE TO DRUGS, LEFT HUMERUS|OSTEONECROSIS DUE TO DRUGS, LEFT HUMERUS
C2901989|T046|M87.121|ICD10CM|OSTEONECROSIS DUE TO DRUGS, RIGHT HUMERUS|OSTEONECROSIS DUE TO DRUGS, RIGHT HUMERUS
C2977004|T047|I82.509|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED DEEP VEINS OF UNSPECIFIED LOWER EXTREMITY|CHRONIC EMBOLISM AND THOMBOS UNSP DEEP VN UNSP LOW EXTRM
C0839948|T047|M86.20|ICD10AM|SUBACUTE OSTEOMYELITIS, UNSPECIFIED SITE|SUBACUTE OSTEOMYELITIS, MULTIPLE SITES
C2838687|T037|S34.129D|ICD10CM|INCOMPLETE LESION OF UNSPECIFIED LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|INCOMPLETE LESION OF UNSP LEVEL OF LUMBAR SPINAL CORD, SUBS
C1829846|T047||ICD10CM|OTHER DISORDERS OF FATTY-ACID OXIDATION
C2838688|T037|S34.129S|ICD10CM|INCOMPLETE LESION OF UNSPECIFIED LEVEL OF LUMBAR SPINAL CORD, SEQUELA|INCOMPLETE LESION OF UNSP LEVEL OF LUM SPINAL CORD, SEQUELA
C2874243|T047|E71.314|ICD10CM|MUSCLE CARNITINE PALMITOYLTRANSFERASE DEFICIENCY|MUSCLE CARNITINE PALMITOYLTRANSFERASE DEFICIENCY
C0220710|T047|E71.311|ICD10CM|MEDIUM CHAIN ACYL COA DEHYDROGENASE DEFICIENCY|MEDIUM CHAIN ACYL COA DEHYDROGENASE DEFICIENCY
C2874239|T047|E71.310|ICD10CM|LONG CHAIN/VERY LONG CHAIN ACYL COA DEHYDROGENASE DEFICIENCY|LCAD
C2874242|T047|E71.313|ICD10CM|GLUTARIC ACIDURIA TYPE II|GLUTARIC ACIDURIA TYPE II C
C0342783|T047|E71.312|ICD10CM|SHORT CHAIN ACYL COA DEHYDROGENASE DEFICIENCY|SCAD
C2879388|T037|T46.0X2A|ICD10CM|POISONING BY CARDIAC-STIMULANT GLYCOSIDES AND DRUGS OF SIMILAR ACTION, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY CARDI-STIM GLYCOS/DRUG SIMLAR ACT, SELF-HARM, INIT
C2833974|T037|S14.135S|ICD10CM|ANTERIOR CORD SYNDROME AT C5 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|ANTERIOR CORD SYNDROME AT C5, SEQUELA
C2887804|T047|K51.30|ICD10CM|ULCERATIVE (CHRONIC) RECTOSIGMOIDITIS WITHOUT COMPLICATIONS|ULCERATIVE (CHRONIC) RECTOSIGMOIDITIS WITHOUT COMPLICATIONS
C2883584|T037|T50.2X2A|ICD10CM|POISONING BY CARBONIC-ANHYDRASE INHIBITORS, BENZOTHIADIAZIDES AND OTHER DIURETICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY CRBNC-ANHYDR INHIBTR,BENZO/OTH DIURETC,SLF-HRM,INIT
C2889084|T047|M02.829|ICD10CM|OTHER REACTIVE ARTHROPATHIES, UNSPECIFIED ELBOW|OTHER REACTIVE ARTHROPATHIES, UNSPECIFIED ELBOW
C2902032|T046|M87.20|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED BONE|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED BONE
C2855997|T037|S68.529S|ICD10CM|PARTIAL TRAUMATIC TRANSPHALANGEAL AMPUTATION OF UNSPECIFIED THUMB, SEQUELA|PARTIAL TRAUMATIC TRNSPHAL AMPUTATION OF THMB, SEQUELA
C2833972|T037|S14.135A|ICD10CM|ANTERIOR CORD SYNDROME AT C5 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|ANTERIOR CORD SYNDROME AT C5, INIT
C2859148|T037|S73.003A|ICD10CM|UNSPECIFIED SUBLUXATION OF UNSPECIFIED HIP, INITIAL ENCOUNTER|UNSPECIFIED SUBLUXATION OF UNSPECIFIED HIP, INIT ENCNTR
C2887649|T047|K27.6|ICD10CM|CHRONIC OR UNSPECIFIED PEPTIC ULCER, SITE UNSPECIFIED, WITH BOTH HEMORRHAGE AND PERFORATION|CHR OR UNSP PEPTIC ULCER, SITE UNSP, W BOTH HEMOR AND PERF
C0840037|T046|M87.28|ICD10AM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, OTHER SITE|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, OTHER SITE
C0494731|T047|K27.5|DMDICD10|CHRONIC OR UNSPECIFIED PEPTIC ULCER, SITE UNSPECIFIED, WITH PERFORATION|ULCUS PEPTICUM, LOKALISATION NICHT NAEHER BEZEICHNET: CHRONISCH ODER NICHT NAEHER BEZEICHNET, MIT PERFORATION
C2887647|T047|K27.2|ICD10CM|ACUTE PEPTIC ULCER, SITE UNSPECIFIED, WITH BOTH HEMORRHAGE AND PERFORATION|ACUTE PEPTIC ULCER, SITE UNSP, W BOTH HEMORRHAGE AND PERF
C0267291|T047|K27.1|DMDICD10|ACUTE PEPTIC ULCER, SITE UNSPECIFIED, WITH PERFORATION|ULCUS PEPTICUM, LOKALISATION NICHT NAEHER BEZEICHNET: AKUT, MIT PERFORATION
C2877173|T037|T38.7X2A|ICD10CM|POISONING BY ANDROGENS AND ANABOLIC CONGENERS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY ANDROGENS AND ANABOLIC CONGENERS, SELF-HARM, INIT
C2887794|T047|K51.018|ICD10CM|ULCERATIVE (CHRONIC) PANCOLITIS WITH OTHER COMPLICATION|ULCERATIVE (CHRONIC) PANCOLITIS WITH OTHER COMPLICATION
C2887795|T047|K51.019|ICD10CM|ULCERATIVE (CHRONIC) PANCOLITIS WITH UNSPECIFIED COMPLICATIONS|ULCERATIVE (CHRONIC) PANCOLITIS WITH UNSP COMPLICATIONS
C2845884|T191|C63.10|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED SPERMATIC CORD|MALIGNANT NEOPLASM OF UNSPECIFIED SPERMATIC CORD
C2845885|T191|C63.11|ICD10CM|MALIGNANT NEOPLASM OF RIGHT SPERMATIC CORD|MALIGNANT NEOPLASM OF RIGHT SPERMATIC CORD
C2845886|T191|C63.12|ICD10CM|MALIGNANT NEOPLASM OF LEFT SPERMATIC CORD|MALIGNANT NEOPLASM OF LEFT SPERMATIC CORD
C2887791|T047|K51.012|ICD10CM|ULCERATIVE (CHRONIC) PANCOLITIS WITH INTESTINAL OBSTRUCTION|ULCERATIVE (CHRONIC) PANCOLITIS WITH INTESTINAL OBSTRUCTION
C2887792|T047|K51.013|ICD10CM|ULCERATIVE (CHRONIC) PANCOLITIS WITH FISTULA|ULCERATIVE (CHRONIC) PANCOLITIS WITH FISTULA
C2887790|T047|K51.011|ICD10CM|ULCERATIVE (CHRONIC) PANCOLITIS WITH RECTAL BLEEDING|ULCERATIVE (CHRONIC) PANCOLITIS WITH RECTAL BLEEDING
C2887793|T047|K51.014|ICD10CM|ULCERATIVE (CHRONIC) PANCOLITIS WITH ABSCESS|ULCERATIVE (CHRONIC) PANCOLITIS WITH ABSCESS
C2835334|T037|S22.050A|ICD10CM|WEDGE COMPRESSION FRACTURE OF T5-T6 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|WEDGE COMPRESSION FRACTURE OF T5-T6 VERTEBRA, INIT
C2885424|T037|T63.082A|ICD10CM|TOXIC EFFECT OF VENOM OF OTHER AFRICAN AND ASIAN SNAKE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFF OF VENOM OF AFRICAN AND ASIAN SNAKE, SLF-HRM, INIT
C2835335|T037|S22.050B|ICD10CM|WEDGE COMPRESSION FRACTURE OF T5-T6 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|WEDGE COMPRSN FRACTURE OF T5-T6 VERTEBRA, INIT FOR OPN FX
C2875023|T047|G04.89|ICD10CM|OTHER MYELITIS|OTHER MYELITIS
C2830376|T033|R40.2212|ICD10CM|COMA SCALE, BEST VERBAL RESPONSE, NONE, AT ARRIVAL TO EMERGENCY DEPARTMENT|COMA SCALE, BEST VERBAL RESPONSE, NONE, EMR
C2830377|T033|R40.2213|ICD10CM|COMA SCALE, BEST VERBAL RESPONSE, NONE, AT HOSPITAL ADMISSION|COMA SCALE, BEST VERBAL RESPONSE, NONE, ADMIT
C2830374|T033|R40.2210|ICD10CM|COMA SCALE, BEST VERBAL RESPONSE, NONE, UNSPECIFIED TIME|COMA SCALE, BEST VERBAL RESPONSE, NONE, UNSPECIFIED TIME
C2830375|T033|R40.2211|ICD10CM|COMA SCALE, BEST VERBAL RESPONSE, NONE, IN THE FIELD [EMT OR AMBULANCE]|COMA SCALE, BEST VERBAL RESPONSE, NONE, IN THE FIELD
C2830378|T033|R40.2214|ICD10CM|COMA SCALE, BEST VERBAL RESPONSE, NONE, 24 HOURS OR MORE AFTER HOSPITAL ADMISSION|COMA SCALE, BEST VERBAL RESPONSE, NONE, 24+HRS
C2890402|T037|T84.010A|ICD10CM|BROKEN INTERNAL RIGHT HIP PROSTHESIS, INITIAL ENCOUNTER|BROKEN INTERNAL RIGHT HIP PROSTHESIS, INITIAL ENCOUNTER
C2890119|T037|T82.595A|ICD10CM|OTHER MECHANICAL COMPLICATION OF UMBRELLA DEVICE, INITIAL ENCOUNTER|MECH COMPL OF UMBRELLA DEVICE, INITIAL ENCOUNTER
C2896597|T046|M80.061A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, RIGHT LOWER LEG, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, R LOW LEG, INIT
C2843318|T037|S48.129S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN UNSPECIFIED SHOULDER AND ELBOW, SEQUELA|PART TRAUM AMP AT LEVEL BETW UNSP SHLDR AND ELBOW, SEQUELA
C2873803|T046|D68.69|ICD10CM|OTHER THROMBOPHILIA|HYPERCOAGULABLE STATES NEC
C2888956|T047|M01.X71|ICD10CM|DIRECT INFECTION OF RIGHT ANKLE AND FOOT IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIR INFCT OF RIGHT ANK/FT IN INFEC/PARASTC DIS CLASSD ELSWHR
C2911418|T033|Z89.441|ICD10CM|ACQUIRED ABSENCE OF RIGHT ANKLE|ACQUIRED ABSENCE OF RIGHT ANKLE
C0085278|T047|D68.61|ICD10CM|ANTIPHOSPHOLIPID SYNDROME|ANTICARDIOLIPIN SYNDROME
C2873802|T047|D68.62|ICD10CM|LUPUS ANTICOAGULANT SYNDROME|PRESENCE OF SYSTEMIC LUPUS ERYTHEMATOSUS [SLE] INHIBITOR
C2911420|T033|Z89.449|ICD10CM|ACQUIRED ABSENCE OF UNSPECIFIED ANKLE|ACQUIRED ABSENCE OF UNSPECIFIED ANKLE
C2837950|T191|C34.10|ICD10CM|MALIGNANT NEOPLASM OF UPPER LOBE, UNSPECIFIED BRONCHUS OR LUNG|MALIGNANT NEOPLASM OF UPPER LOBE, UNSP BRONCHUS OR LUNG
C2837951|T191|C34.11|ICD10CM|MALIGNANT NEOPLASM OF UPPER LOBE, RIGHT BRONCHUS OR LUNG|MALIGNANT NEOPLASM OF UPPER LOBE, RIGHT BRONCHUS OR LUNG
C2837952|T191|C34.12|ICD10CM|MALIGNANT NEOPLASM OF UPPER LOBE, LEFT BRONCHUS OR LUNG|MALIGNANT NEOPLASM OF UPPER LOBE, LEFT BRONCHUS OR LUNG
C2977723|T037|S02.69XA|ICD10CM|FRACTURE OF MANDIBLE OF OTHER SPECIFIED SITE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF MANDIBLE OF OTH SITE, INIT FOR CLOS FX
C2901256|T046|M84.552A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, LEFT FEMUR, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, LEFT FEMUR, INIT
C2890103|T037|T82.591A|ICD10CM|OTHER MECHANICAL COMPLICATION OF SURGICALLY CREATED ARTERIOVENOUS SHUNT, INITIAL ENCOUNTER|MECH COMPL OF SURGICALLY CREATED ARTERIOVENOUS SHUNT, INIT
C2901524|T046|M84.663A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, RIGHT FIBULA, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, RIGHT FIBULA, INIT
C2902170|T046|M87.879|ICD10CM|OTHER OSTEONECROSIS, UNSPECIFIED TOE(S)|OTHER OSTEONECROSIS, UNSPECIFIED TOE(S)
C2902169|T046|M87.878|ICD10CM|OTHER OSTEONECROSIS, LEFT TOE(S)|OTHER OSTEONECROSIS, LEFT TOE(S)
C2977728|T037|S02.69XS|ICD10CM|FRACTURE OF MANDIBLE OF OTHER SPECIFIED SITE, SEQUELA|FRACTURE OF MANDIBLE OF OTHER SPECIFIED SITE, SEQUELA
C2888958|T047|M01.X79|ICD10CM|DIRECT INFECTION OF UNSPECIFIED ANKLE AND FOOT IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIR INFCT OF UNSP ANK/FT IN INFEC/PARASTC DIS CLASSD ELSWHR
C2902162|T046|M87.871|ICD10CM|OTHER OSTEONECROSIS, RIGHT ANKLE|OTHER OSTEONECROSIS, RIGHT ANKLE
C2902164|T046|M87.873|ICD10CM|OTHER OSTEONECROSIS, UNSPECIFIED ANKLE|OTHER OSTEONECROSIS, UNSPECIFIED ANKLE
C2902163|T046|M87.872|ICD10CM|OTHER OSTEONECROSIS, LEFT ANKLE|OTHER OSTEONECROSIS, LEFT ANKLE
C2902166|T046|M87.875|ICD10CM|OTHER OSTEONECROSIS, LEFT FOOT|OTHER OSTEONECROSIS, LEFT FOOT
C2902165|T046|M87.874|ICD10CM|OTHER OSTEONECROSIS, RIGHT FOOT|OTHER OSTEONECROSIS, RIGHT FOOT
C2902168|T046|M87.877|ICD10CM|OTHER OSTEONECROSIS, RIGHT TOE(S)|OTHER OSTEONECROSIS, RIGHT TOE(S)
C2902167|T046|M87.876|ICD10CM|OTHER OSTEONECROSIS, UNSPECIFIED FOOT|OTHER OSTEONECROSIS, UNSPECIFIED FOOT
C2901110|T046|M84.478A|ICD10CM|PATHOLOGICAL FRACTURE, LEFT TOE(S), INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, LEFT TOE(S), INIT ENCNTR FOR FRACTURE
C2882155|T033|I22.9|ICD10CM|SUBSEQUENT ST ELEVATION (STEMI) MYOCARDIAL INFARCTION OF UNSPECIFIED SITE|SUBSEQUENT STEMI OF UNSP SITE
C2882152|T033|I22.8|ICD10CM|SUBSEQUENT ST ELEVATION (STEMI) MYOCARDIAL INFARCTION OF OTHER SITES|SUBSEQUENT STEMI OF SITES
C2882141|T033|I22.2|ICD10CM|SUBSEQUENT NON-ST ELEVATION (NSTEMI) MYOCARDIAL INFARCTION|SUBSEQUENT NON-ST ELEVATION (NSTEMI) MYOCARDIAL INFARCTION
C3839202|T047|I22.1|ICD10CM|SUBSEQUENT ST ELEVATION (STEMI) MYOCARDIAL INFARCTION OF INFERIOR WALL|SUBSEQUENT STEMI OF INFERIOR WALL
C2882131|T047|I22.0|ICD10CM|SUBSEQUENT ST ELEVATION (STEMI) MYOCARDIAL INFARCTION OF ANTERIOR WALL|SUBSEQUENT STEMI OF ANTERIOR WALL
C2838646|T037|S34.112D|ICD10CM|COMPLETE LESION OF L2 LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION OF L2 LEVEL OF LUMBAR SPINAL CORD, SUBS
C2838645|T037|S34.112A|ICD10CM|COMPLETE LESION OF L2 LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION OF L2 LEVEL OF LUMBAR SPINAL CORD, INIT
C2837987|T191|C43.12|ICD10CM|MALIGNANT MELANOMA OF LEFT EYELID, INCLUDING CANTHUS|MALIGNANT MELANOMA OF LEFT EYELID, INCLUDING CANTHUS
C2837985|T191|C43.10|ICD10CM|MALIGNANT MELANOMA OF UNSPECIFIED EYELID, INCLUDING CANTHUS|MALIGNANT MELANOMA OF UNSPECIFIED EYELID, INCLUDING CANTHUS
C2837986|T191|C43.11|ICD10CM|MALIGNANT MELANOMA OF RIGHT EYELID, INCLUDING CANTHUS|MALIGNANT MELANOMA OF RIGHT EYELID, INCLUDING CANTHUS
C2884530|T037|T56.4X2S|ICD10CM|TOXIC EFFECT OF COPPER AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF COPPER AND ITS COMPOUNDS, SELF-HARM, SEQUELA
C2880001|T037|T48.292S|ICD10CM|POISONING BY OTHER DRUGS ACTING ON MUSCLES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH DRUGS ACTING ON MUSCLES, SELF-HARM, SEQUELA
C2879517|T037|T46.5X2A|ICD10CM|POISONING BY OTHER ANTIHYPERTENSIVE DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH ANTIHYPERTENSIVE DRUGS, SELF-HARM, INIT
C2884528|T037|T56.4X2A|ICD10CM|TOXIC EFFECT OF COPPER AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF COPPER AND ITS COMPOUNDS, SELF-HARM, INIT
C3543852|T047|R53.2|ICD10CM|FUNCTIONAL QUADRIPLEGIA|FUNCTIONAL QUADRIPLEGIA
C2879999|T037|T48.292A|ICD10CM|POISONING BY OTHER DRUGS ACTING ON MUSCLES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH DRUGS ACTING ON MUSCLES, SELF-HARM, INIT
C2874490|T048|F12.250|ICD10CM|CANNABIS DEPENDENCE WITH PSYCHOTIC DISORDER WITH DELUSIONS|CANNABIS DEPENDENCE WITH PSYCHOTIC DISORDER WITH DELUSIONS
C2874491|T048|F12.251|ICD10CM|CANNABIS DEPENDENCE WITH PSYCHOTIC DISORDER WITH HALLUCINATIONS|CANNABIS DEPENDENCE W PSYCHOTIC DISORDER WITH HALLUCINATIONS
C2889391|T047|M06.02|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, UNSPECIFIED ELBOW|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, ELBOW
C2874492|T048|F12.259|ICD10CM|CANNABIS DEPENDENCE WITH PSYCHOTIC DISORDER, UNSPECIFIED|CANNABIS DEPENDENCE WITH PSYCHOTIC DISORDER, UNSPECIFIED
C2889392|T047|M06.021|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, RIGHT ELBOW|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, RIGHT ELBOW
C2889393|T047|M06.022|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, LEFT ELBOW|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, LEFT ELBOW
C0496818|T191|C54.0|DMDICD10|MALIGNANT NEOPLASM OF ISTHMUS UTERI|BOESARTIGE NEUBILDUNG: ISTHMUS UTERI
C0007103|T191|C54.1|DMDICD10|MALIGNANT NEOPLASM OF ENDOMETRIUM|BOESARTIGE NEUBILDUNG: ENDOMETRIUM
C0496820|T191|C54.2|DMDICD10|MALIGNANT NEOPLASM OF MYOMETRIUM|BOESARTIGE NEUBILDUNG: MYOMETRIUM
C0496821|T191|C54.3|DMDICD10|MALIGNANT NEOPLASM OF FUNDUS UTERI|BOESARTIGE NEUBILDUNG: FUNDUS UTERI
C0348907|T191|C54.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF CORPUS UTERI|BOESARTIGE NEUBILDUNG: CORPUS UTERI, MEHRERE TEILBEREICHE UEBERLAPPEND
C0153574|T191|C54.9|DMDICD10|MALIGNANT NEOPLASM OF CORPUS UTERI, UNSPECIFIED|BOESARTIGE NEUBILDUNG: CORPUS UTERI, NICHT NAEHER BEZEICHNET
C2835450|T037|S22.081B|ICD10CM|STABLE BURST FRACTURE OF T11-T12 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|STABLE BURST FRACTURE OF T11-T12 VERTEBRA, INIT FOR OPN FX
C2835449|T037|S22.081A|ICD10CM|STABLE BURST FRACTURE OF T11-T12 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|STABLE BURST FRACTURE OF T11-T12 VERTEBRA, INIT FOR CLOS FX
C2882849|T047|I70.468|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, OTHER EXTREMITY|ATHSCL AUTOL VEIN BYPASS OF THE EXTRM W GANGRENE, OTH EXTRM
C2882850|T047|I70.469|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, UNSPECIFIED EXTREMITY|ATHSCL AUTOL VEIN BYPASS OF THE EXTRM W GANGRENE, UNSP EXTRM
C2882846|T047|I70.461|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, RIGHT LEG|ATHSCL AUTOL VEIN BYPASS OF THE EXTRM W GANGRENE, RIGHT LEG
C2882847|T047|I70.462|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, LEFT LEG|ATHSCL AUTOL VEIN BYPASS OF THE EXTRM W GANGRENE, LEFT LEG
C2882848|T047|I70.463|ICD10CM|ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, BILATERAL LEGS|ATHSCL AUTOL VEIN BYPASS OF THE EXTRM W GANGRENE, BI LEGS
C0920028|T191|C95.92|ICD10CM|LEUKEMIA, UNSPECIFIED, IN RELAPSE|LEUKEMIA, UNSPECIFIED, IN RELAPSE
C0686584|T191||ICD10AM|LEUKEMIA, UNSPECIFIED, IN REMISSION
C2861647|T191|C95.90|ICD10CM|LEUKEMIA, UNSPECIFIED NOT HAVING ACHIEVED REMISSION|LEUKEMIA, UNSPECIFIED NOT HAVING ACHIEVED REMISSION
C2876944|T037|T37.8X2A|ICD10CM|POISONING BY OTHER SPECIFIED SYSTEMIC ANTI-INFECTIVES AND ANTIPARASITICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY OTH SYSTEMIC ANTI-INFECT/PARASIT, SELF-HARM, INIT
C4270590|T046|T85.734A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO IMPLANTED ELECTRONIC NEUROSTIMULATOR, GENERATOR, INITIAL ENCOUNTER|I/I REACT D/T IMPLNT ELEC NSTIM, GENERATOR, INIT
C2883507|T037|T49.92XA|ICD10CM|POISONING BY UNSPECIFIED TOPICAL AGENT, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY UNSP TOPICAL AGENT, INTENTIONAL SELF-HARM, INIT
C2832148|T037|S06.323A|ICD10CM|CONTUSION AND LACERATION OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|CONTUS/LAC LEFT CEREBRUM W LOC OF 1-5 HRS 59 MIN, INIT
C2883509|T037|T49.92XS|ICD10CM|POISONING BY UNSPECIFIED TOPICAL AGENT, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY UNSP TOPICAL AGENT, SELF-HARM, SEQUELA
C2882662|T046|I69.939|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING UNSPECIFIED SIDE|MONOPLG UPR LMB FOL UNSP CEREBVASC DISEASE AFF UNSP SIDE
C0347509|T191|D33.9|DMDICD10|BENIGN NEOPLASM OF CENTRAL NERVOUS SYSTEM, UNSPECIFIED|GUTARTIGE NEUBILDUNG: ZENTRALNERVENSYSTEM, NICHT NAEHER BEZEICHNET
C0348419|T191|D33.7|DMDICD10|BENIGN NEOPLASM OF OTHER SPECIFIED PARTS OF CENTRAL NERVOUS SYSTEM|GUTARTIGE NEUBILDUNG: SONSTIGE NAEHER BEZEICHNETE TEILE DES ZENTRALNERVENSYSTEMS
C0154034|T191|D33.4|DMDICD10|BENIGN NEOPLASM OF SPINAL CORD|GUTARTIGE NEUBILDUNG: RUECKENMARK
C2882660|T046|I69.933|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING RIGHT NON-DOMINANT SIDE|MONOPLG UPR LMB FOL UNSP CEREBVASC DIS AFF RIGHT NONDOM SIDE
C0496899|T191|D33.2|DMDICD10|BENIGN NEOPLASM OF BRAIN, UNSPECIFIED|GUTARTIGE NEUBILDUNG: GEHIRN, NICHT NAEHER BEZEICHNET
C2869557|T191|D33.3|ICD10CM|BENIGN NEOPLASM OF CRANIAL NERVES|BENIGN NEOPLASM OF OLFACTORY BULB
C0686393|T191|D33.0|ICD10CM|BENIGN NEOPLASM OF BRAIN, SUPRATENTORIAL|BENIGN NEOPLASM OF CEREBRAL VENTRICLE
C2869556|T191|D33.1|ICD10CM|BENIGN NEOPLASM OF BRAIN, INFRATENTORIAL|BENIGN NEOPLASM OF FOURTH VENTRICLE
C0494228|T047|D57.1|DMDICD10|SICKLE-CELL DISEASE WITHOUT CRISIS|SICHELZELLENANAEMIE OHNE KRISEN
C2905818|T037|X83.8XXD|ICD10CM|INTENTIONAL SELF-HARM BY OTHER SPECIFIED MEANS, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY OTHER SPECIFIED MEANS, SUBS ENCNTR
C2832268|T037|S06.351S|ICD10CM|TRAUMATIC HEMORRHAGE OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|TRAUM HEMOR L CEREB W LOC OF 30 MINUTES OR LESS, SEQUELA
C2831399|T037|S02.0XXS|ICD10CM|FRACTURE OF VAULT OF SKULL, SEQUELA|FRACTURE OF VAULT OF SKULL, SEQUELA
C0037054|T047|D57.3|DMDICD10|SICKLE-CELL TRAIT|SICHELZELLEN-ERBANLAGE
C2832266|T037|S06.351A|ICD10CM|TRAUMATIC HEMORRHAGE OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|TRAUM HEMOR LEFT CEREBRUM W LOC OF 30 MINUTES OR LESS, INIT
C2831395|T037|S02.0XXB|ICD10CM|FRACTURE OF VAULT OF SKULL, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF VAULT OF SKULL, INIT ENCNTR FOR OPEN FRACTURE
C2831394|T037|S02.0XXA|ICD10CM|FRACTURE OF VAULT OF SKULL, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF VAULT OF SKULL, INIT ENCNTR FOR CLOSED FRACTURE
C2889649|T047|M08.971|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, RIGHT ANKLE AND FOOT|JUVENILE ARTHRITIS, UNSPECIFIED, RIGHT ANKLE AND FOOT
C2889650|T047|M08.972|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, LEFT ANKLE AND FOOT|JUVENILE ARTHRITIS, UNSPECIFIED, LEFT ANKLE AND FOOT
C2889651|T047|M08.979|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, UNSPECIFIED ANKLE AND FOOT|JUVENILE ARTHRITIS, UNSPECIFIED, UNSPECIFIED ANKLE AND FOOT
C4269291|T037|S02.11BS|ICD10CM|TYPE I OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, SEQUELA|TYPE I OCCIPITAL CONDYLE FRACTURE, LEFT SIDE, SEQUELA
C2887167|T047|I82.C29|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED INTERNAL JUGULAR VEIN|CHRONIC EMBOLISM AND THOMBOS UNSP INTERNAL JUGULAR VEIN
C2890759|T037|T84.328A|ICD10CM|DISPLACEMENT OF OTHER BONE DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|DISPLACEMENT OF OTH BONE DEVICES, IMPLANTS AND GRAFTS, INIT
C2887165|T047|I82.C22|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF LEFT INTERNAL JUGULAR VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF L INT JUGULAR VEIN
C2887166|T047|I82.C23|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF INTERNAL JUGULAR VEIN, BILATERAL|CHRONIC EMBOLISM AND THOMBOS OF INT JUGULAR VEIN, BILATERAL
C2887164|T047|I82.C21|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF RIGHT INTERNAL JUGULAR VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF R INT JUGULAR VEIN
C0494231|T046|D59.2|DMDICD10|DRUG-INDUCED NONAUTOIMMUNE HEMOLYTIC ANEMIA|ARZNEIMITTELINDUZIERTE NICHT-AUTOIMMUNHAEMOLYTISCHE ANAEMIE
C0019061|T047|D59.3|DMDICD10|HEMOLYTIC-UREMIC SYNDROME|HAEMOLYTISCH-URAEMISCHES SYNDROM
C0391817|T046|D59.0|DMDICD10|DRUG-INDUCED AUTOIMMUNE HEMOLYTIC ANEMIA|ARZNEIMITTELINDUZIERTE AUTOIMMUNHAEMOLYTISCHE ANAEMIE
C2873775|T047|D59.1|ICD10CM|OTHER AUTOIMMUNE HEMOLYTIC ANEMIAS|AUTOIMMUNE HEMOLYTIC DISEASE (COLD TYPE) (WARM TYPE)
C0494233|T047|D59.6|DMDICD10|HEMOGLOBINURIA DUE TO HEMOLYSIS FROM OTHER EXTERNAL CAUSES|HAEMOGLOBINURIE DURCH HAEMOLYSE INFOLGE SONSTIGER AEUSSERER URSACHEN
C0021051|T047|D84.9|DMDICD10|IMMUNODEFICIENCY, UNSPECIFIED|IMMUNDEFEKT, NICHT NAEHER BEZEICHNET
C1321858|T047|D59.4|ICD10CM|OTHER NONAUTOIMMUNE HEMOLYTIC ANEMIAS|MECHANICAL HEMOLYTIC ANEMIA
C0024790|T047|D59.5|DMDICD10|PAROXYSMAL NOCTURNAL HEMOGLOBINURIA [MARCHIAFAVA-MICHELI]|PAROXYSMALE NAECHTLICHE HAEMOGLOBINURIE [MARCHIAFAVA-MICHELI]
C2878816|T037|T44.3X2A|ICD10CM|POISONING BY OTHER PARASYMPATHOLYTICS [ANTICHOLINERGICS AND ANTIMUSCARINICS] AND SPASMOLYTICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY OTH PARASYMPATH AND SPASMOLYTICS, SELF-HARM, INIT
C0477309|T047|D59.8|DMDICD10|OTHER ACQUIRED HEMOLYTIC ANEMIAS|SONSTIGE ERWORBENE HAEMOLYTISCHE ANAEMIEN
C0271904|T047||ICD10CM|ACQUIRED HEMOLYTIC ANEMIA, UNSPECIFIED
C0451699|T047|D84.0|DMDICD10|LYMPHOCYTE FUNCTION ANTIGEN-1 [LFA-1] DEFECT|LYMPHOZYTENFUNKTION-ANTIGEN-1[LFA-1]-DEFEKT
C2873848|T047|D84.1|ICD10CM|DEFECTS IN THE COMPLEMENT SYSTEM|C1 ESTERASE INHIBITOR [C1-INH] DEFICIENCY
C4268663|T047|K86.89|ICD10CM|OTHER SPECIFIED DISEASES OF PANCREAS|PANCREATIC NECROSIS NOS, UNRELATED TO ACUTE PANCREATITIS
C0267963|T047|K86.81|ICD10CM|EXOCRINE PANCREATIC INSUFFICIENCY|EXOCRINE PANCREATIC INSUFFICIENCY
C2878818|T037|T44.3X2S|ICD10CM|POISONING BY OTHER PARASYMPATHOLYTICS [ANTICHOLINERGICS AND ANTIMUSCARINICS] AND SPASMOLYTICS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY OTH PARASYMPATH AND SPASMOLYTICS, SLF-HRM, SEQUELA
C4269298|T037|S02.11CS|ICD10CM|TYPE II OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, SEQUELA|TYPE II OCCIPITAL CONDYLE FRACTURE, RIGHT SIDE, SEQUELA
C2874004|T047|E09.622|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH OTHER SKIN ULCER|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS W OTH SKIN ULCER
C2910364|T019|Q92.62|ICD10CM|MARKER CHROMOSOMES IN ABNORMAL INDIVIDUAL|MARKER CHROMOSOMES IN ABNORMAL INDIVIDUAL
C2874002|T047|E09.620|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH DIABETIC DERMATITIS|DRUG/CHEM DIABETES MELLITUS W DIABETIC DERMATITIS
C2874003|T047|E09.621|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH FOOT ULCER|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH FOOT ULCER
C0153024|T047||ICD10CM|POSTHERPETIC TRIGEMINAL NEURALGIA
C2874005|T047|E09.628|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH OTHER SKIN COMPLICATIONS|DRUG/CHEM DIABETES MELLITUS W OTH SKIN COMPLICATIONS
C2837832|T037|S32.312A|ICD10CM|DISPLACED AVULSION FRACTURE OF LEFT ILIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED AVULSION FRACTURE OF LEFT ILIUM, INIT FOR CLOS FX
C2837833|T037|S32.312B|ICD10CM|DISPLACED AVULSION FRACTURE OF LEFT ILIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISPLACED AVULSION FRACTURE OF LEFT ILIUM, INIT FOR OPN FX
C0837587|T047|M06.20|ICD10AM|RHEUMATOID BURSITIS, UNSPECIFIED SITE|RHEUMATOID BURSITIS, MULTIPLE SITES
C2889438|T047||ICD10CM|RHEUMATOID BURSITIS, VERTEBRAE
C0837587|T047|M06.29|ICD10CM|RHEUMATOID BURSITIS, MULTIPLE SITES|RHEUMATOID BURSITIS, MULTIPLE SITES
C0362053|T048||ICD10CM|OTHER DISSOCIATIVE AND CONVERSION DISORDERS
C0026773|T048||ICD10CM|DISSOCIATIVE IDENTITY DISORDER
C2900493|T047|B02.24|ICD10CM|POSTHERPETIC MYELITIS|POSTHERPETIC MYELITIS
C2833562|T037|S12.551B|ICD10CM|OTHER TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH TRAUM NONDISP SPONDYLOLYSIS OF SIXTH CERVCAL VERT, 7THB
C4270503|T046|T85.191A|ICD10CM|OTHER MECHANICAL COMPLICATION OF IMPLANTED ELECTRONIC NEUROSTIMULATOR OF PERIPHERAL NERVE ELECTRODE (LEAD), INITIAL ENCOUNTER|MECH COMPL OF IMPLNT ELEC NSTIM OF PRPH NRV LEAD, INIT
C2883636|T037|T50.4X2S|ICD10CM|POISONING BY DRUGS AFFECTING URIC ACID METABOLISM, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY DRUGS AFF URIC ACID METAB, SELF-HARM, SEQUELA
C2842116|T191|C50.521|ICD10CM|MALIGNANT NEOPLASM OF LOWER-OUTER QUADRANT OF RIGHT MALE BREAST|MALIG NEOPLASM OF LOWER-OUTER QUADRANT OF RIGHT MALE BREAST
C2832262|T037|S06.350A|ICD10CM|TRAUMATIC HEMORRHAGE OF LEFT CEREBRUM WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|TRAUM HEMOR LEFT CEREBRUM W/O LOSS OF CONSCIOUSNESS, INIT
C2883634|T037|T50.4X2A|ICD10CM|POISONING BY DRUGS AFFECTING URIC ACID METABOLISM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY DRUGS AFF URIC ACID METAB, SELF-HARM, INIT
C2903164|T046|N99.518|ICD10CM|OTHER CYSTOSTOMY COMPLICATION|OTHER CYSTOSTOMY COMPLICATION
C2842117|T191|C50.522|ICD10CM|MALIGNANT NEOPLASM OF LOWER-OUTER QUADRANT OF LEFT MALE BREAST|MALIG NEOPLASM OF LOWER-OUTER QUADRANT OF LEFT MALE BREAST
C2903162|T046|N99.510|ICD10CM|CYSTOSTOMY HEMORRHAGE|CYSTOSTOMY HEMORRHAGE
C2903163|T046|N99.511|ICD10CM|CYSTOSTOMY INFECTION|CYSTOSTOMY INFECTION
C1397892|T046|N99.512|ICD10CM|CYSTOSTOMY MALFUNCTION|CYSTOSTOMY MALFUNCTION
C2858339|T037|S72.411B|ICD10CM|DISPLACED UNSPECIFIED CONDYLE FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL UNSP CONDYLE FX LOW END R FEMR, 7THB
C2882735|T047|I70.262|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES WITH GANGRENE, LEFT LEG|ATHSCL NATIVE ARTERIES OF EXTREMITIES W GANGRENE, LEFT LEG
C2882736|T047|I70.263|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES WITH GANGRENE, BILATERAL LEGS|ATHSCL NATIVE ARTERIES OF EXTRM W GANGRENE, BILATERAL LEGS
C2889136|T047|M05.112|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT SHOULDER|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF L SHOULDER
C2882734|T047|I70.261|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES WITH GANGRENE, RIGHT LEG|ATHSCL NATIVE ARTERIES OF EXTREMITIES W GANGRENE, RIGHT LEG
C2900911|T046|M84.431A|ICD10CM|PATHOLOGICAL FRACTURE, RIGHT ULNA, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, RIGHT ULNA, INIT ENCNTR FOR FRACTURE
C2889137|T047|M05.119|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER|RHEU LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP SHOULDER
C2882737|T047|I70.268|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES WITH GANGRENE, OTHER EXTREMITY|ATHSCL NATIVE ARTERIES OF EXTRM W GANGRENE, OTH EXTREMITY
C2882738|T047|I70.269|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF EXTREMITIES WITH GANGRENE, UNSPECIFIED EXTREMITY|ATHSCL NATIVE ARTERIES OF EXTRM W GANGRENE, UNSP EXTREMITY
C2860038|T037|S78.921S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF RIGHT HIP AND THIGH, LEVEL UNSPECIFIED, SEQUELA|PARTIAL TRAUM AMP OF R HIP AND THIGH, LEVEL UNSP, SEQUELA
C2883709|T037|T50.7X2A|ICD10CM|POISONING BY ANALEPTICS AND OPIOID RECEPTOR ANTAGONISTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY ANALEPTICS AND OPIOID RECEPTOR ANTAG, SLF-HRM, INIT
C4268620|T047|K55.031|ICD10CM|FOCAL (SEGMENTAL) ACUTE (REVERSIBLE) ISCHEMIA OF LARGE INTESTINE|FOCAL (SEGMENTAL) ACUTE ISCHEMIA OF LARGE INTESTINE
C4270810|T047|K55.032|ICD10CM|DIFFUSE ACUTE (REVERSIBLE) ISCHEMIA OF LARGE INTESTINE|DIFFUSE ACUTE (REVERSIBLE) ISCHEMIA OF LARGE INTESTINE
C4268621|T047|K55.039|ICD10CM|ACUTE (REVERSIBLE) ISCHEMIA OF LARGE INTESTINE, EXTENT UNSPECIFIED|ACUTE ISCHEMIA OF LARGE INTESTINE, EXTENT UNSPECIFIED
C2832198|T037|S06.335A|ICD10CM|CONTUSION AND LACERATION OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, INITIAL ENCOUNTER|CONTUS/LAC CEREB, W LOC >24 HR W RET CONSC LEV, INIT
C2890264|T037|T83.121A|ICD10CM|DISPLACEMENT OF IMPLANTED URINARY SPHINCTER, INITIAL ENCOUNTER|DISPLACEMENT OF IMPLANTED URINARY SPHINCTER, INIT
C2832200|T037|S06.335S|ICD10CM|CONTUSION AND LACERATION OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, SEQUELA|CONTUS/LAC CEREB, W LOC >24 HR W RET CONSC LEV, SEQUELA
C3264136|T033|Z89.511|ICD10CM|ACQUIRED ABSENCE OF RIGHT LEG BELOW KNEE|ACQUIRED ABSENCE OF RIGHT LEG BELOW KNEE
C2874697|T048|F16.229|ICD10CM|HALLUCINOGEN DEPENDENCE WITH INTOXICATION, UNSPECIFIED|HALLUCINOGEN DEPENDENCE WITH INTOXICATION, UNSPECIFIED
C2874696|T048|F16.221|ICD10CM|HALLUCINOGEN DEPENDENCE WITH INTOXICATION WITH DELIRIUM|HALLUCINOGEN DEPENDENCE WITH INTOXICATION WITH DELIRIUM
C2874695|T048||ICD10CM|HALLUCINOGEN DEPENDENCE WITH INTOXICATION, UNCOMPLICATED
C2843295|T037|S48.111A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN RIGHT SHOULDER AND ELBOW, INITIAL ENCOUNTER|COMPLETE TRAUM AMP AT LEVEL BETW R SHOULDER AND ELBOW, INIT
C2859044|T037|S72.8X2A|ICD10CM|OTHER FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF LEFT FEMUR, INIT ENCNTR FOR CLOSED FRACTURE
C2858851|T037|S72.461A|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPL SUPRCNDL FX W INTRCNDL EXTN LOWER END OF R FEMUR, INIT
C2865568|T037|S88.911A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT LOWER LEG, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF R LOW LEG, LEVEL UNSP, INIT
C2865569|T037|S88.911D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT LOWER LEG, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF R LOW LEG, LEVEL UNSP, SUBS
C2843297|T037|S48.111S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN RIGHT SHOULDER AND ELBOW, SEQUELA|COMPLETE TRAUM AMP AT LEVEL BETW R SHLDR AND ELBOW, SEQUELA
C0153368|T191|C04.9|DMDICD10|MALIGNANT NEOPLASM OF FLOOR OF MOUTH, UNSPECIFIED|BOESARTIGE NEUBILDUNG: MUNDBODEN, NICHT NAEHER BEZEICHNET
C0349046|T191|C04.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF FLOOR OF MOUTH|BOESARTIGE NEUBILDUNG: MUNDBODEN, MEHRERE TEILBEREICHE UEBERLAPPEND
C2858594|T037|S72.434B|ICD10CM|NONDISPLACED FRACTURE OF MEDIAL CONDYLE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF MED CONDYLE OF R FEMR, 7THB
C0496758|T191|C04.1|DMDICD10|MALIGNANT NEOPLASM OF LATERAL FLOOR OF MOUTH|BOESARTIGE NEUBILDUNG: SEITLICHER TEIL DES MUNDBODENS
C2833836|T191|C04.0|ICD10CM|MALIGNANT NEOPLASM OF ANTERIOR FLOOR OF MOUTH|MALIGNANT NEOPLASM OF ANTERIOR TO THE PREMOLAR-CANINE JUNCTION
C2835781|T037|S24.112D|ICD10CM|COMPLETE LESION AT T2-T6 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION AT T2-T6 LEVEL OF THORACIC SPINAL CORD, SUBS
C2834037|T037|S14.152D|ICD10CM|OTHER INCOMPLETE LESION AT C2 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|OTH INCOMPLETE LESION AT C2, SUBS
C2833420|T037|S12.350A|ICD10CM|OTHER TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH TRAUM DISPL SPONDYLOLYSIS OF FOURTH CERVCAL VERT, INIT
C2858010|T037|S72.346A|ICD10CM|NONDISPLACED SPIRAL FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED SPIRAL FRACTURE OF SHAFT OF UNSP FEMUR, INIT
C2858011|T037|S72.346B|ICD10CM|NONDISPLACED SPIRAL FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP SPIRAL FX SHAFT OF UNSP FEMR, 7THB
C2835780|T037|S24.112A|ICD10CM|COMPLETE LESION AT T2-T6 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION AT T2-T6 LEVEL OF THORACIC SPINAL CORD, INIT
C2891275|T037||ICD10CM|CARDIAC ALLOGRAFT VASCULOPATHY
C2891274|T037|T86.298|ICD10CM|OTHER COMPLICATIONS OF HEART TRANSPLANT|OTHER COMPLICATIONS OF HEART TRANSPLANT
C2835782|T037|S24.112S|ICD10CM|COMPLETE LESION AT T2-T6 LEVEL OF THORACIC SPINAL CORD, SEQUELA|COMPLETE LESION AT T2-T6, SEQUELA
C2889691|T037|T81.592A|ICD10CM|OTHER COMPLICATIONS OF FOREIGN BODY ACCIDENTALLY LEFT IN BODY FOLLOWING KIDNEY DIALYSIS, INITIAL ENCOUNTER|OTH COMP OF FB ACC LEFT IN BODY FOL KIDNEY DIALYSIS, INIT
C2901828|T047|M86.239|ICD10CM|SUBACUTE OSTEOMYELITIS, UNSPECIFIED RADIUS AND ULNA|SUBACUTE OSTEOMYELITIS, UNSPECIFIED RADIUS AND ULNA
C0477408|T047|G73.3|DMDICD10|MYASTHENIC SYNDROMES IN OTHER DISEASES CLASSIFIED ELSEWHERE|MYASTHENIESYNDROME BEI SONSTIGEN ANDERENORTS KLASSIFIZIERTEN KRANKHEITEN
C3161081|T047||ICD10CM|LAMBERT-EATON SYNDROME IN NEOPLASTIC DISEASE
C2838208|T037|S32.455B|ICD10CM|NONDISPLACED TRANSVERSE FRACTURE OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP TRANSVERSE FX LEFT ACETABULUM, INIT FOR OPN FX
C2875322|T047|G73.7|ICD10CM|MYOPATHY IN DISEASES CLASSIFIED ELSEWHERE|MYOPATHY IN DISEASES CLASSIFIED ELSEWHERE
C2874179|T033|E16.3|ICD10CM|INCREASED SECRETION OF GLUCAGON|HYPERPLASIA OF PANCREATIC ENDOCRINE CELLS WITH GLUCAGON EXCESS
C2874181|T047|E16.4|ICD10CM|INCREASED SECRETION OF GASTRIN|INCREASED SECRETION OF GASTRIN
C2838672|T037|S34.122S|ICD10CM|INCOMPLETE LESION OF L2 LEVEL OF LUMBAR SPINAL CORD, SEQUELA|INCOMPLETE LESION OF L2 LEVEL OF LUMBAR SPINAL CORD, SEQUELA
C2874185|T047|E16.8|ICD10CM|OTHER SPECIFIED DISORDERS OF PANCREATIC INTERNAL SECRETION|INCREASED SECRETION FROM ENDOCRINE PANCREAS OF VASOACTIVE-INTESTINAL POLYPEPTIDE
C1263961|T047|E16.9|DMDICD10|DISORDER OF PANCREATIC INTERNAL SECRETION, UNSPECIFIED|STOERUNG DER INNEREN SEKRETION DES PANKREAS, NICHT NAEHER BEZEICHNET
C2837581|T037|S32.039A|ICD10CM|UNSPECIFIED FRACTURE OF THIRD LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF THIRD LUMBAR VERTEBRA, INIT FOR CLOS FX
C2865516|T037|S88.011A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT KNEE LEVEL, RIGHT LOWER LEG, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION AT KNEE LEVEL, R LOW LEG, INIT
C2905703|T037|X74.02XA|ICD10CM|INTENTIONAL SELF-HARM BY PAINTBALL GUN, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY PAINTBALL GUN, INITIAL ENCOUNTER
C2889072|T047|M02.369|ICD10CM|REITER'S DISEASE, UNSPECIFIED KNEE|REITER'S DISEASE, UNSPECIFIED KNEE
C0036421|T047|M34|DMDICD10|SYSTEMIC SCLEROSIS, UNSPECIFIED|SYSTEMISCHE SKLEROSE
C2889071|T047|M02.362|ICD10CM|REITER'S DISEASE, LEFT KNEE|REITER'S DISEASE, LEFT KNEE
C2889070|T047|M02.361|ICD10CM|REITER'S DISEASE, RIGHT KNEE|REITER'S DISEASE, RIGHT KNEE
C0036421|T047|M34|DMDICD10|PROGRESSIVE SYSTEMIC SCLEROSIS|SYSTEMISCHE SKLEROSE
C2895195|T047|M34.1|ICD10CM|CR(E)ST SYNDROME|COMBINATION OF CALCINOSIS, RAYNAUD'S PHENOMENON, ESOPHAGEAL DYSFUNCTION, SCLERODACTYLY, TELANGIECTASIA
C0451842|T037|M34.2|DMDICD10|SYSTEMIC SCLEROSIS INDUCED BY DRUG AND CHEMICAL|SYSTEMISCHE SKLEROSE, DURCH ARZNEIMITTEL ODER CHEMISCHE SUBSTANZEN INDUZIERT
C2901827|T047|M86.232|ICD10CM|SUBACUTE OSTEOMYELITIS, LEFT RADIUS AND ULNA|SUBACUTE OSTEOMYELITIS, LEFT RADIUS AND ULNA
C2901154|T046|M84.519A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, UNSPECIFIED SHOULDER, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, UNSP SHOULDER, INIT
C2874820|T048|F19.23|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH WITHDRAWAL, UNSPECIFIED|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH WITHDRAWAL
C0162283|T047|N25.1|DMDICD10|NEPHROGENIC DIABETES INSIPIDUS|RENALER DIABETES INSIPIDUS
C1527410|T047|N25.0|ICD10CM|RENAL OSTEODYSTROPHY|RENAL RICKETS
C2890690|T037|T84.199A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTERNAL FIXATION DEVICE OF UNSPECIFIED BONE OF LIMB, INITIAL ENCOUNTER|MECH COMPL OF INT FIX OF UNSP BONE OF LIMB, INIT
C0342204|T047|E02|DMDICD10|SUBCLINICAL IODINE-DEFICIENCY HYPOTHYROIDISM|SUBKLINISCHE JODMANGEL-HYPOTHYREOSE
C2860014|T037|S78.122A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN LEFT HIP AND KNEE, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP AT LEVEL BETW LEFT HIP AND KNEE, INIT
C2887062|T047|A32.7|ICD10CM|LISTERIAL SEPSIS|LISTERIAL SEPSIS
C2860015|T037|S78.122D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN LEFT HIP AND KNEE, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMP AT LEVEL BETW LEFT HIP AND KNEE, SUBS
C2890775|T037|T84.410A|ICD10CM|BREAKDOWN (MECHANICAL) OF MUSCLE AND TENDON GRAFT, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF MUSCLE AND TENDON GRAFT, INIT
C2887176|T047|I83.008|ICD10CM|VARICOSE VEINS OF UNSPECIFIED LOWER EXTREMITY WITH ULCER OTHER PART OF LOWER LEG|VARICOS VN UNSP LOW EXTRM W ULCER OTH PART OF LOWER LEG
C2887177|T047|I83.009|ICD10CM|VARICOSE VEINS OF UNSPECIFIED LOWER EXTREMITY WITH ULCER OF UNSPECIFIED SITE|VARICOSE VEINS OF UNSP LOWER EXTREMITY W ULCER OF UNSP SITE
C4236995|T048|F90.2|ICD10CM|ATTENTION-DEFICIT HYPERACTIVITY DISORDER, COMBINED TYPE|ATTENTION-DEFICIT/HYPERACTIVITY DISORDER, COMBINED PRESENTATION
C4236996|T048|F90.1|ICD10CM|ATTENTION-DEFICIT HYPERACTIVITY DISORDER, PREDOMINANTLY HYPERACTIVE TYPE|ATTENTION-DEFICIT/HYPERACTIVITY DISORDER, PREDOMINANTLY HYPERACTIVE IMPULSIVE PRESENTATION
C4236997|T048|F90.0|ICD10CM|ATTENTION-DEFICIT HYPERACTIVITY DISORDER, PREDOMINANTLY INATTENTIVE TYPE|ATTENTION-DEFICIT/HYPERACTIVITY DISORDER, PREDOMINANTLY INATTENTIVE PRESENTATION
C2887169|T047|I83.001|ICD10CM|VARICOSE VEINS OF UNSPECIFIED LOWER EXTREMITY WITH ULCER OF THIGH|VARICOSE VEINS OF UNSP LOWER EXTREMITY WITH ULCER OF THIGH
C2887170|T047|I83.002|ICD10CM|VARICOSE VEINS OF UNSPECIFIED LOWER EXTREMITY WITH ULCER OF CALF|VARICOSE VEINS OF UNSP LOWER EXTREMITY WITH ULCER OF CALF
C2887171|T047|I83.003|ICD10CM|VARICOSE VEINS OF UNSPECIFIED LOWER EXTREMITY WITH ULCER OF ANKLE|VARICOSE VEINS OF UNSP LOWER EXTREMITY WITH ULCER OF ANKLE
C2887173|T047|I83.004|ICD10CM|VARICOSE VEINS OF UNSPECIFIED LOWER EXTREMITY WITH ULCER OF HEEL AND MIDFOOT|VARICOS VN UNSP LOWER EXTREMITY W ULCER OF HEEL AND MIDFOOT
C2887175|T047|I83.005|ICD10CM|VARICOSE VEINS OF UNSPECIFIED LOWER EXTREMITY WITH ULCER OTHER PART OF FOOT|VARICOS VN UNSP LOWER EXTREMITY W ULCER OTH PART OF FOOT
C2875001|T048|F90.9|ICD10CM|ATTENTION-DEFICIT HYPERACTIVITY DISORDER, UNSPECIFIED TYPE|ATTENTION-DEFICIT HYPERACTIVITY DISORDER, UNSPECIFIED TYPE
C2874999|T048|F90.8|ICD10CM|ATTENTION-DEFICIT HYPERACTIVITY DISORDER, OTHER TYPE|ATTENTION-DEFICIT HYPERACTIVITY DISORDER, OTHER TYPE
C4268281|T048|F18.27|ICD10CM|INHALANT DEPENDENCE WITH INHALANT-INDUCED DEMENTIA|INHALANT USE DISORDER, SEVERE, WITH INHALANT INDUCED MAJOR NEUROCOGNITIVE DISORDER
C4268279|T048|F18.24|ICD10CM|INHALANT DEPENDENCE WITH INHALANT-INDUCED MOOD DISORDER|INHALANT USE DISORDER, SEVERE, WITH INHALANT INDUCED DEPRESSIVE DISORDER
C4237148|T048|F18.20|ICD10CM|INHALANT DEPENDENCE, UNCOMPLICATED|INHALANT USE DISORDER, SEVERE
C4509105|T048|F18.21|ICD10CM|INHALANT DEPENDENCE, IN REMISSION|INHALANT USE DISORDER, SEVERE, IN SUSTAINED REMISSION
C2838279|T037|S32.473A|ICD10CM|DISPLACED FRACTURE OF MEDIAL WALL OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF MEDIAL WALL OF UNSP ACETABULUM, INIT FOR CLOS FX
C2874771|T048|F18.29|ICD10CM|INHALANT DEPENDENCE WITH UNSPECIFIED INHALANT-INDUCED DISORDER|INHALANT DEPENDENCE WITH UNSP INHALANT-INDUCED DISORDER
C0348494|T047|E78.4|DMDICD10|OTHER HYPERLIPIDEMIA|SONSTIGE HYPERLIPIDAEMIEN
C0020473|T047|E78.5|DMDICD10|HYPERLIPIDEMIA, UNSPECIFIED|HYPERLIPIDAEMIE, NICHT NAEHER BEZEICHNET
C3165209|T047||ICD10CM|LIPOPROTEIN DEFICIENCY
C2893642|T047|M12.049|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], UNSPECIFIED HAND|CHRONIC POSTRHEUMATIC ARTHROPATHY, UNSPECIFIED HAND
C2874288|T033|E78.1|ICD10CM|PURE HYPERGLYCERIDEMIA|ELEVATED FASTING TRIGLYCERIDES
C2874289|T033|E78.2|ICD10CM|MIXED HYPERLIPIDEMIA|HYPERCHOLESTEREMIA WITH ENDOGENOUS HYPERGLYCERIDEMIA
C0795956|T047|E78.3|ICD10CM|HYPERCHYLOMICRONEMIA|CHYLOMICRON RETENTION DISEASE
C2893641|T047|M12.042|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], LEFT HAND|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], LEFT HAND
C2893640|T047|M12.041|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], RIGHT HAND|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], RIGHT HAND
C0494345|T047|E78.9|DMDICD10|DISORDER OF LIPOPROTEIN METABOLISM, UNSPECIFIED|STOERUNG DES LIPOPROTEINSTOFFWECHSELS, NICHT NAEHER BEZEICHNET
C2888562|T047|L89.619|ICD10CM|PRESSURE ULCER OF RIGHT HEEL, UNSPECIFIED STAGE|PRESSURE ULCER OF RIGHT HEEL, UNSPECIFIED STAGE
C2977724|T037|S02.69XB|ICD10CM|FRACTURE OF MANDIBLE OF OTHER SPECIFIED SITE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF MANDIBLE OF OTH SITE, INIT FOR OPN FX
C2833561|T037|S12.551A|ICD10CM|OTHER TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH TRAUM NONDISP SPONDYLOLYSIS OF SIXTH CERVCAL VERT, INIT
C3263955|T048||ICD10CM|OTHER PERVASIVE DEVELOPMENTAL DISORDERS
C0524528|T048|F84|DMDICD10|PERVASIVE DEVELOPMENTAL DISORDER, UNSPECIFIED|TIEFGREIFENDE ENTWICKLUNGSSTOERUNGEN
C2902871|T046|N02.6|ICD10CM|RECURRENT AND PERSISTENT HEMATURIA WITH DENSE DEPOSIT DISEASE|RECURRENT AND PERSISTENT HEMATURIA WITH MEMBRANOPROLIFERATIVE GLOMERULONEPHRITIS, TYPE 2
C0035372|T047|F84.2|DMDICD10|RETT'S SYNDROME|RETT-SYNDROM
C0349329|T048|F84.3|DMDICD10|OTHER CHILDHOOD DISINTEGRATIVE DISORDER|ANDERE DESINTEGRATIVE STOERUNG DES KINDESALTERS
C2603372|T048|F84.0|ICD10CM|AUTISTIC DISORDER|INFANTILE PSYCHOSIS
C1306579|T047||ICD10CM|ASPERGER'S SYNDROME
C2882452|T047|I69.031|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING RIGHT DOMINANT SIDE|MONOPLG UPR LMB FOL NTRM SUBARACH HEMOR AFF RIGHT DOM SIDE
C2882454|T047|I69.033|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING RIGHT NON-DOMINANT SIDE|MONOPLG UPR LMB FOL NTRM SUBARACH HEMOR AFF R NONDOM SIDE
C2882453|T047|I69.032|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING LEFT DOMINANT SIDE|MONOPLG UPR LMB FOL NTRM SUBARACH HEMOR AFF LEFT DOM SIDE
C2882455|T047|I69.034|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING LEFT NON-DOMINANT SIDE|MONOPLG UPR LMB FOL NTRM SUBARACH HEMOR AFF LEFT NONDOM SIDE
C2882456|T047|I69.039|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING NONTRAUMATIC SUBARACHNOID HEMORRHAGE AFFECTING UNSPECIFIED SIDE|MONOPLG UPR LMB FOLLOWING NTRM SUBARACH HEMOR AFF UNSP SIDE
C2859046|T037|S72.8X2C|ICD10CM|OTHER FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|OTH FRACTURE OF LEFT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2859045|T037|S72.8X2B|ICD10CM|OTHER FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|OTH FRACTURE OF LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C2905704|T037|X74.02XD|ICD10CM|INTENTIONAL SELF-HARM BY PAINTBALL GUN, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY PAINTBALL GUN, SUBSEQUENT ENCOUNTER
C2896559|T046|M80.042A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, LEFT HAND, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, LEFT HAND, INIT
C2884867|T037|T59.2X2S|ICD10CM|TOXIC EFFECT OF FORMALDEHYDE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF FORMALDEHYDE, INTENTIONAL SELF-HARM, SEQUELA
C2888547|T047||ICD10CM|PRESSURE ULCER OF RIGHT HEEL, UNSTAGEABLE
C2888550|T047|L89.611|ICD10CM|PRESSURE ULCER OF RIGHT HEEL, STAGE 1|PRESSURE ULCER OF RIGHT HEEL, STAGE 1
C2888553|T047|L89.612|ICD10CM|PRESSURE ULCER OF RIGHT HEEL, STAGE 2|PRESSURE ULCER OF RIGHT HEEL, STAGE 2
C2888556|T047|L89.613|ICD10CM|PRESSURE ULCER OF RIGHT HEEL, STAGE 3|PRESSURE ULCER OF RIGHT HEEL, STAGE 3
C2888559|T047|L89.614|ICD10CM|PRESSURE ULCER OF RIGHT HEEL, STAGE 4|PRESSURE ULCER OF RIGHT HEEL, STAGE 4
C2838280|T037|S32.473B|ICD10CM|DISPLACED FRACTURE OF MEDIAL WALL OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISP FX OF MEDIAL WALL OF UNSP ACETABULUM, INIT FOR OPN FX
C0525045|T048|F39|DMDICD10|UNSPECIFIED MOOD [AFFECTIVE] DISORDER|NICHT NAEHER BEZEICHNETE AFFEKTIVE STOERUNG
C2884865|T037|T59.2X2A|ICD10CM|TOXIC EFFECT OF FORMALDEHYDE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF FORMALDEHYDE, INTENTIONAL SELF-HARM, INIT
C2883062|T047|I80.203|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF UNSPECIFIED DEEP VESSELS OF LOWER EXTREMITIES, BILATERAL|PHLBTS AND THOMBOPHLB OF UNSP DEEP VESSELS OF LOW EXTRM, BI
C2883061|T047|I80.202|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF UNSPECIFIED DEEP VESSELS OF LEFT LOWER EXTREMITY|PHLBTS AND THOMBOPHLB OF UNSP DEEP VESSELS OF L LOW EXTREM
C2883060|T047|I80.201|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF UNSPECIFIED DEEP VESSELS OF RIGHT LOWER EXTREMITY|PHLBTS AND THOMBOPHLB OF UNSP DEEP VESSELS OF R LOW EXTREM
C2837460|T037|S32.002B|ICD10CM|UNSTABLE BURST FRACTURE OF UNSPECIFIED LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSTABLE BURST FX UNSP LUM VERTEBRA, INIT FOR OPN FX
C2883063|T047|I80.209|ICD10CM|PHLEBITIS AND THROMBOPHLEBITIS OF UNSPECIFIED DEEP VESSELS OF UNSPECIFIED LOWER EXTREMITY|PHLBTS AND THOMBOPHLB OF UNSP DEEP VESSELS OF UNSP LOW EXTRM
C2349263|T191|C90.12|ICD10CM|PLASMA CELL LEUKEMIA IN RELAPSE|PLASMA CELL LEUKEMIA IN RELAPSE
C2854077|T191||ICD10CM|PLASMA CELL LEUKEMIA NOT HAVING ACHIEVED REMISSION
C0153871|T191||ICD10AMAE|PLASMA CELL LEUKEMIA IN REMISSION
C2890195|T037|T82.898A|ICD10CM|OTHER SPECIFIED COMPLICATION OF VASCULAR PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|OTH COMPLICATION OF VASCULAR PROSTH DEV/GRFT, INIT
C0837077|T047|E13.36|ICD10AM|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC CATARACT|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC CATARACT
C2901356|T046|M84.58XA|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, OTHER SPECIFIED SITE, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, OTH SITE, INIT
C2835819|T037|S24.141D|ICD10CM|BROWN-SEQUARD SYNDROME AT T1 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|BROWN-SEQUARD SYNDROME AT T1, SUBS
C4268283|T048|F18.288|ICD10CM|INHALANT DEPENDENCE WITH OTHER INHALANT-INDUCED DISORDER|INHALANT USE DISORDER, SEVERE, WITH INHALANT-INDUCED MILD NEUROCOGNITIVE DISORDER
C2876225|T037|T32.88|ICD10CM|CORROSIONS INVOLVING 80-89% OF BODY SURFACE WITH 80-89% THIRD DEGREE CORROSION|CORROS 80-89% OF BODY SURFACE W 80-89% THIRD DEGREE CORROS
C2876219|T037|T32.82|ICD10CM|CORROSIONS INVOLVING 80-89% OF BODY SURFACE WITH 20-29% THIRD DEGREE CORROSION|CORROS 80-89% OF BODY SURFACE W 20-29% THIRD DEGREE CORROS
C2876220|T037|T32.83|ICD10CM|CORROSIONS INVOLVING 80-89% OF BODY SURFACE WITH 30-39% THIRD DEGREE CORROSION|CORROS 80-89% OF BODY SURFACE W 30-39% THIRD DEGREE CORROS
C2876218|T037|T32.81|ICD10CM|CORROSIONS INVOLVING 80-89% OF BODY SURFACE WITH 10-19% THIRD DEGREE CORROSION|CORROS 80-89% OF BODY SURFACE W 10-19% THIRD DEGREE CORROS
C2876223|T037|T32.86|ICD10CM|CORROSIONS INVOLVING 80-89% OF BODY SURFACE WITH 60-69% THIRD DEGREE CORROSION|CORROS 80-89% OF BODY SURFACE W 60-69% THIRD DEGREE CORROS
C2876224|T037|T32.87|ICD10CM|CORROSIONS INVOLVING 80-89% OF BODY SURFACE WITH 70-79% THIRD DEGREE CORROSION|CORROS 80-89% OF BODY SURFACE W 70-79% THIRD DEGREE CORROS
C2876221|T037|T32.84|ICD10CM|CORROSIONS INVOLVING 80-89% OF BODY SURFACE WITH 40-49% THIRD DEGREE CORROSION|CORROS 80-89% OF BODY SURFACE W 40-49% THIRD DEGREE CORROS
C2876222|T037|T32.85|ICD10CM|CORROSIONS INVOLVING 80-89% OF BODY SURFACE WITH 50-59% THIRD DEGREE CORROSION|CORROS 80-89% OF BODY SURFACE W 50-59% THIRD DEGREE CORROS
C2885443|T037|T63.092S|ICD10CM|TOXIC EFFECT OF VENOM OF OTHER SNAKE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF SNAKE, SELF-HARM, SEQUELA
C2885441|T037|T63.092A|ICD10CM|TOXIC EFFECT OF VENOM OF OTHER SNAKE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF SNAKE, INTENTIONAL SELF-HARM, INIT
C3264406|T046||ICD10CM|ACUTE POSTPROCEDURAL RESPIRATORY FAILURE
C3264407|T046||ICD10CM|ACUTE AND CHRONIC POSTPROCEDURAL RESPIRATORY FAILURE
C2874107|T047|E11.59|ICD10CM|TYPE 2 DIABETES MELLITUS WITH OTHER CIRCULATORY COMPLICATIONS|TYPE 2 DIABETES MELLITUS WITH OTH CIRCULATORY COMPLICATIONS
C0265316|T047|Q85.9|DMDICD10|PHAKOMATOSIS, UNSPECIFIED|PHAKOMATOSE, NICHT NAEHER BEZEICHNET
C2876135|T037|T31.32|ICD10CM|BURNS INVOLVING 30-39% OF BODY SURFACE WITH 20-29% THIRD DEGREE BURNS|BURNS OF 30-39% OF BODY SURFACE W 20-29% THIRD DEGREE BURNS
C2876136|T037|T31.33|ICD10CM|BURNS INVOLVING 30-39% OF BODY SURFACE WITH 30-39% THIRD DEGREE BURNS|BURNS OF 30-39% OF BODY SURFACE W 30-39% THIRD DEGREE BURNS
C0349219|T048|F33.0|DMDICD10|MAJOR DEPRESSIVE DISORDER, RECURRENT, MILD|REZIDIVIERENDE DEPRESSIVE STOERUNG, GEGENWAERTIG LEICHTE EPISODE
C0154411|T048|F33.1|DMDICD10|MAJOR DEPRESSIVE DISORDER, RECURRENT, MODERATE|REZIDIVIERENDE DEPRESSIVE STOERUNG, GEGENWAERTIG MITTELGRADIGE EPISODE
C0154412|T048|F33.2|DMDICD10|MAJOR DEPRESSIVE DISORDER, RECURRENT SEVERE WITHOUT PSYCHOTIC FEATURES|REZIDIVIERENDE DEPRESSIVE STOERUNG, GEGENWAERTIG SCHWERE EPISODE OHNE PSYCHOTISCHE SYMPTOME
C2874931|T048|F33.3|ICD10CM|MAJOR DEPRESSIVE DISORDER, RECURRENT, SEVERE WITH PSYCHOTIC SYMPTOMS|MAJOR DEPRESSV DISORDER, RECURRENT, SEVERE W PSYCH SYMPTOMS
C2874104|T047|E11.51|ICD10CM|TYPE 2 DIABETES MELLITUS WITH DIABETIC PERIPHERAL ANGIOPATHY WITHOUT GANGRENE|TYPE 2 DIABETES W DIABETIC PERIPHERAL ANGIOPATH W/O GANGRENE
C0041341|T191|Q85.1|DMDICD10|TUBEROUS SCLEROSIS|TUBEROESE (HIRN-) SKLEROSE
C2874106|T047|E11.52|ICD10CM|TYPE 2 DIABETES MELLITUS WITH DIABETIC PERIPHERAL ANGIOPATHY WITH GANGRENE|TYPE 2 DIABETES W DIABETIC PERIPHERAL ANGIOPATHY W GANGRENE
C2874934|T048|F33.8|ICD10CM|OTHER RECURRENT DEPRESSIVE DISORDERS|RECURRENT BRIEF DEPRESSIVE EPISODES
C0349218|T048|F33|DMDICD10|MAJOR DEPRESSIVE DISORDER, RECURRENT, UNSPECIFIED|REZIDIVIERENDE DEPRESSIVE STOERUNG
C2901770|T047|M86.011|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, RIGHT SHOULDER|ACUTE HEMATOGENOUS OSTEOMYELITIS, RIGHT SHOULDER
C2901771|T047|M86.012|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, LEFT SHOULDER|ACUTE HEMATOGENOUS OSTEOMYELITIS, LEFT SHOULDER
C4270411|T046|T83.724A|ICD10CM|EXPOSURE OF IMPLANTED URETERAL BULKING AGENT INTO URETER, INITIAL ENCOUNTER|EXPOSURE OF IMPLNT URETERAL BULKING AGENT INTO URETER, INIT
C2901772|T047|M86.019|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED SHOULDER|ACUTE HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED SHOULDER
C2349314|T191||ICD10CM|MALIGNANT CARCINOID TUMOR OF THE DUODENUM
C2349315|T191||ICD10CM|MALIGNANT CARCINOID TUMOR OF THE JEJUNUM
C2349316|T191||ICD10CM|MALIGNANT CARCINOID TUMOR OF THE ILEUM
C2349313|T191|C7A.019|ICD10CM|MALIGNANT CARCINOID TUMOR OF THE SMALL INTESTINE, UNSPECIFIED PORTION|MALIGNANT CARCINOID TUMOR OF THE SM INT, UNSP PORTION
C3264204|T047|H40.1233|ICD10CM|LOW-TENSION GLAUCOMA, BILATERAL, SEVERE STAGE|LOW-TENSION GLAUCOMA, BILATERAL, SEVERE STAGE
C2842111|T191|C50.429|ICD10CM|MALIGNANT NEOPLASM OF UPPER-OUTER QUADRANT OF UNSPECIFIED MALE BREAST|MALIG NEOPLASM OF UPPER-OUTER QUADRANT OF UNSP MALE BREAST
C3264202|T047|H40.1231|ICD10CM|LOW-TENSION GLAUCOMA, BILATERAL, MILD STAGE|LOW-TENSION GLAUCOMA, BILATERAL, MILD STAGE
C3264201|T047|H40.1230|ICD10CM|LOW-TENSION GLAUCOMA, BILATERAL, STAGE UNSPECIFIED|LOW-TENSION GLAUCOMA, BILATERAL, STAGE UNSPECIFIED
C3264205|T047|H40.1234|ICD10CM|LOW-TENSION GLAUCOMA, BILATERAL, INDETERMINATE STAGE|LOW-TENSION GLAUCOMA, BILATERAL, INDETERMINATE STAGE
C2842109|T191|C50.421|ICD10CM|MALIGNANT NEOPLASM OF UPPER-OUTER QUADRANT OF RIGHT MALE BREAST|MALIG NEOPLASM OF UPPER-OUTER QUADRANT OF RIGHT MALE BREAST
C2842110|T191|C50.422|ICD10CM|MALIGNANT NEOPLASM OF UPPER-OUTER QUADRANT OF LEFT MALE BREAST|MALIG NEOPLASM OF UPPER-OUTER QUADRANT OF LEFT MALE BREAST
C2835820|T037|S24.141S|ICD10CM|BROWN-SEQUARD SYNDROME AT T1 LEVEL OF THORACIC SPINAL CORD, SEQUELA|BROWN-SEQUARD SYNDROME AT T1, SEQUELA
C2884318|T037|T53.7X2A|ICD10CM|TOXIC EFFECT OF OTHER HALOGEN DERIVATIVES OF AROMATIC HYDROCARBONS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFF OF HALGN DERIV OF AROMATIC HYDROCRB, SLF-HRM, INIT
C2349335|T191|C7A.1|ICD10CM|MALIGNANT POORLY DIFFERENTIATED NEUROENDOCRINE TUMORS|MALIGNANT POORLY DIFFERENTIATED NEUROENDOCRINE TUMORS
C2845977|T191|C7A.8|ICD10CM|OTHER MALIGNANT NEUROENDOCRINE TUMORS|OTHER MALIGNANT NEUROENDOCRINE TUMORS
C2884320|T037|T53.7X2S|ICD10CM|TOXIC EFFECT OF OTHER HALOGEN DERIVATIVES OF AROMATIC HYDROCARBONS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFF OF HALGN DERIV OF AROMATIC HYDROCRB, SLF-HRM, SQLA
C2882435|T047|I66.22|ICD10CM|OCCLUSION AND STENOSIS OF LEFT POSTERIOR CEREBRAL ARTERY|OCCLUSION AND STENOSIS OF LEFT POSTERIOR CEREBRAL ARTERY
C2882436|T047|I66.23|ICD10CM|OCCLUSION AND STENOSIS OF BILATERAL POSTERIOR CEREBRAL ARTERIES|OCCLUSION AND STENOSIS OF BI POSTERIOR CEREBRAL ARTERIES
C2882434|T047|I66.21|ICD10CM|OCCLUSION AND STENOSIS OF RIGHT POSTERIOR CEREBRAL ARTERY|OCCLUSION AND STENOSIS OF RIGHT POSTERIOR CEREBRAL ARTERY
C2888712|T047|L97.424|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT HEEL AND MIDFOOT WITH NECROSIS OF BONE|NON-PRS CHRONIC ULCER OF LEFT HEEL AND MIDFOOT W NECROS BONE
C2874150|T047|E13.39|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH OTHER DIABETIC OPHTHALMIC COMPLICATION|OTH DIABETES MELLITUS W OTH DIABETIC OPHTHALMIC COMPLICATION
C4509309|T047|L97.426|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT HEEL AND MIDFOOT WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OF L HEEL/MIDFT W BNE INVL W/O EVD OF NECR
C2874800|T048|F19.15|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE ABUSE WITH PSYCHOACTIVE SUBSTANCE-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|OTHER PSYCHOACTIVE SUBSTANCE ABUSE WITH PSYCHOACTIVE SUBSTANCE-INDUCED PSYCHOTIC DISORDER
C2888710|T047|L97.422|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT HEEL AND MIDFOOT WITH FAT LAYER EXPOSED|NON-PRS CHR ULCER OF LEFT HEEL AND MIDFOOT W FAT LAYER EXPOS
C2882437|T047|I66.29|ICD10CM|OCCLUSION AND STENOSIS OF UNSPECIFIED POSTERIOR CEREBRAL ARTERY|OCCLUSION AND STENOSIS OF UNSP POSTERIOR CEREBRAL ARTERY
C4268075|T047|E11.3299|ICD10CM|TYPE 2 DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|TYPE 2 DIAB WITH MILD NONP RTNOP WITHOUT MACULAR EDEMA, UNSP
C0839976|T047|M86.48|ICD10AM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, OTHER SITE|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, OTHER SITE
C0839968|T047|M86.49|ICD10CM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, MULTIPLE SITES|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, MULTIPLE SITES
C2883128|T047|I82.529|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED ILIAC VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF UNSPECIFIED ILIAC VEIN
C2889204|T047|M05.321|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT ELBOW|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF R ELBOW
C4268072|T047|E11.3291|ICD10CM|TYPE 2 DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|TYPE 2 DIAB WITH MILD NONP RTNOP WITHOUT MCLR EDEMA, R EYE
C4268073|T047|E11.3292|ICD10CM|TYPE 2 DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|TYPE 2 DIAB WITH MILD NONP RTNOP WITHOUT MCLR EDEMA, L EYE
C4268074|T047|E11.3293|ICD10CM|TYPE 2 DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|TYPE 2 DIAB WITH MILD NONP RTNOP WITHOUT MACULAR EDEMA, BI
C2883125|T047|I82.521|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF RIGHT ILIAC VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF RIGHT ILIAC VEIN
C2883126|T047|I82.522|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF LEFT ILIAC VEIN|CHRONIC EMBOLISM AND THROMBOSIS OF LEFT ILIAC VEIN
C2883127|T047|I82.523|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF ILIAC VEIN, BILATERAL|CHRONIC EMBOLISM AND THROMBOSIS OF ILIAC VEIN, BILATERAL
C2890291|T037|T83.198A|ICD10CM|OTHER MECHANICAL COMPLICATION OF OTHER URINARY DEVICES AND IMPLANTS, INITIAL ENCOUNTER|MECH COMPL OF OTH URINARY DEVICES AND IMPLANTS, INIT ENCNTR
C0004775|T047||ICD10CM|BARTTER'S SYNDROME
C0864795|T047|A66.6|ICD10CM|BONE AND JOINT LESIONS OF YAWS|YAWS GUMMATOUS OSTEITIS OR PERIOSTITIS
C0348460|T047|E26.89|ICD10CM|OTHER HYPERALDOSTERONISM|OTHER HYPERALDOSTERONISM
C0031572|T048|F40.10|ICD10CM|SOCIAL PHOBIA, UNSPECIFIED|SOCIAL PHOBIA, UNSPECIFIED
C0270587|T048||ICD10CM|SOCIAL PHOBIA, GENERALIZED
C2832637|T037|S06.891S|ICD10CM|OTHER SPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|INTCRAN INJ W LOC OF 30 MINUTES OR LESS, SEQUELA
C0840009|T046|M87.09|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF BONE, MULTIPLE SITES|IDIOPATHIC ASEPTIC NECROSIS OF BONE, MULTIPLE SITES
C0840017|T046|M87.08|ICD10AM|IDIOPATHIC ASEPTIC NECROSIS OF BONE, OTHER SITE|IDIOPATHIC ASEPTIC NECROSIS OF BONE, OTHER SITE
C2833981|T037|S14.137D|ICD10CM|ANTERIOR CORD SYNDROME AT C7 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|ANTERIOR CORD SYNDROME AT C7, SUBS
C2889310|T047|M05.641|ICD10CM|RHEUMATOID ARTHRITIS OF RIGHT HAND WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF RIGHT HAND W INVOLV OF ORGANS AND SYSTEMS
C0151620|T047|I67.4|DMDICD10|HYPERTENSIVE ENCEPHALOPATHY|HYPERTENSIVE ENZEPHALOPATHIE
C2349435|T047|G43.111|ICD10CM|MIGRAINE WITH AURA, INTRACTABLE, WITH STATUS MIGRAINOSUS|MIGRAINE WITH AURA, INTRACTABLE, WITH STATUS MIGRAINOSUS
C2882442|T046||ICD10CM|NONPYOGENIC THROMBOSIS OF INTRACRANIAL VENOUS SYSTEM
C0494615|T047|I67.7|DMDICD10|CEREBRAL ARTERITIS, NOT ELSEWHERE CLASSIFIED|ZEREBRALE ARTERIITIS, ANDERENORTS NICHT KLASSIFIZIERT
C0348838|T020|I67.0|DMDICD10|DISSECTION OF CEREBRAL ARTERIES, NONRUPTURED|DISSEKTION INTRAKRANIELLER ARTERIEN, NICHTRUPTURIERT
C2882441|T047|I67.2|ICD10CM|CEREBRAL ATHEROSCLEROSIS|ATHEROMA OF CEREBRAL AND PRECEREBRAL ARTERIES
C0494613|T046|I67.3|DMDICD10|PROGRESSIVE VASCULAR LEUKOENCEPHALOPATHY|PROGRESSIVE SUBKORTIKALE VASKULAERE ENZEPHALOPATHIE
C2349433|T047|G43.119|ICD10CM|MIGRAINE WITH AURA, INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|MIGRAINE WITH AURA, INTRACTABLE, WITHOUT STATUS MIGRAINOSUS
C0007820|T047|I67.9|DMDICD10|CEREBROVASCULAR DISEASE, UNSPECIFIED|ZEREBROVASKULAERE KRANKHEIT, NICHT NAEHER BEZEICHNET
C2833547|T037|S12.54XB|ICD10CM|TYPE III TRAUMATIC SPONDYLOLISTHESIS OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE III TRAUM SPONDYLOLYSIS OF SIXTH CERVCAL VERT, 7THB
C2874594|T048|F14.229|ICD10CM|COCAINE DEPENDENCE WITH INTOXICATION, UNSPECIFIED|COCAINE DEPENDENCE WITH INTOXICATION, UNSPECIFIED
C2833546|T037|S12.54XA|ICD10CM|TYPE III TRAUMATIC SPONDYLOLISTHESIS OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE III TRAUM SPONDYLOLYSIS OF SIXTH CERVCAL VERTEBRA, INIT
C2877254|T037|T38.892S|ICD10CM|POISONING BY OTHER HORMONES AND SYNTHETIC SUBSTITUTES, INTENTIONAL SELF-HARM, SEQUELA|POISN BY OTH HORMONES AND SYNTHETIC SUB, SELF-HARM, SEQUELA
C2890910|T037|T84.84XA|ICD10CM|PAIN DUE TO INTERNAL ORTHOPEDIC PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|PAIN DUE TO INTERNAL ORTHOPEDIC PROSTH DEV/GRFT, INIT
C0152964|T047|A40.9|DMDICD10|STREPTOCOCCAL SEPSIS, UNSPECIFIED|SEPSIS DURCH STREPTOKOKKEN, NICHT NAEHER BEZEICHNET
C2887085|T047|A40.8|ICD10CM|OTHER STREPTOCOCCAL SEPSIS|OTHER STREPTOCOCCAL SEPSIS
C2887084|T047|A40.3|ICD10CM|SEPSIS DUE TO STREPTOCOCCUS PNEUMONIAE|SEPSIS DUE TO STREPTOCOCCUS PNEUMONIAE
C2887083|T047|A40.1|ICD10CM|SEPSIS DUE TO STREPTOCOCCUS, GROUP B|SEPSIS DUE TO STREPTOCOCCUS, GROUP B
C2887082|T047|A40.0|ICD10CM|SEPSIS DUE TO STREPTOCOCCUS, GROUP A|SEPSIS DUE TO STREPTOCOCCUS, GROUP A
C2911410|T033|Z89.421|ICD10CM|ACQUIRED ABSENCE OF OTHER RIGHT TOE(S)|ACQUIRED ABSENCE OF OTHER RIGHT TOE(S)
C2911411|T033|Z89.422|ICD10CM|ACQUIRED ABSENCE OF OTHER LEFT TOE(S)|ACQUIRED ABSENCE OF OTHER LEFT TOE(S)
C0477350|T047|G12.8|DMDICD10|OTHER SPINAL MUSCULAR ATROPHIES AND RELATED SYNDROMES|SONSTIGE SPINALE MUSKELATROPHIEN UND VERWANDTE SYNDROME
C0026847|T047|G12.9|DMDICD10|SPINAL MUSCULAR ATROPHY, UNSPECIFIED|SPINALE MUSKELATROPHIE, NICHT NAEHER BEZEICHNET
C2911412|T033|Z89.429|ICD10CM|ACQUIRED ABSENCE OF OTHER TOE(S), UNSPECIFIED SIDE|ACQUIRED ABSENCE OF OTHER TOE(S), UNSPECIFIED SIDE
C0043116|T047|G12.0|DMDICD10|INFANTILE SPINAL MUSCULAR ATROPHY, TYPE I [WERDNIG-HOFFMAN]|INFANTILE SPINALE MUSKELATROPHIE, TYP I [TYP WERDNIG-HOFFMANN]
C2875051|T047|G12.1|ICD10CM|OTHER INHERITED SPINAL MUSCULAR ATROPHY|JUVENILE FORM, TYPE III SPINAL MUSCULAR ATROPHY [KUGELBERG-WELANDER]
C2901510|T047|M84.661A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, RIGHT TIBIA, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, RIGHT TIBIA, INIT
C2902152|T046|M87.852|ICD10CM|OTHER OSTEONECROSIS, LEFT FEMUR|OTHER OSTEONECROSIS, LEFT FEMUR
C2902151|T046|M87.851|ICD10CM|OTHER OSTEONECROSIS, RIGHT FEMUR|OTHER OSTEONECROSIS, RIGHT FEMUR
C2902150|T046|M87.850|ICD10CM|OTHER OSTEONECROSIS, PELVIS|OTHER OSTEONECROSIS, PELVIS
C2856027|T037|S68.616S|ICD10CM|COMPLETE TRAUMATIC TRANSPHALANGEAL AMPUTATION OF RIGHT LITTLE FINGER, SEQUELA|COMPLETE TRAUMATIC TRNSPHAL AMP OF R LITTLE FINGER, SEQUELA
C2902153|T046|M87.859|ICD10CM|OTHER OSTEONECROSIS, UNSPECIFIED FEMUR|OTHER OSTEONECROSIS, UNSPECIFIED FEMUR
C1387794|T047||ICD10CM|ANGINA PECTORIS WITH DOCUMENTED SPASM
C2882088|T047|I20.0|ICD10CM|UNSTABLE ANGINA|WORSENING EFFORT ANGINA
C2885609|T037|T63.412A|ICD10CM|TOXIC EFFECT OF VENOM OF CENTIPEDES AND VENOMOUS MILLIPEDES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF CENTIPEDE/MILLIPEDE, SLF-HRM, INIT
C0002962|T184|I20.9|DMDICD10|ANGINA PECTORIS, UNSPECIFIED|ANGINA PECTORIS, NICHT NAEHER BEZEICHNET
C2976973|T047|I20.8|ICD10CM|OTHER FORMS OF ANGINA PECTORIS|CORONARY SLOW FLOW SYNDROME
C2889640|T047|M08.949|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, UNSPECIFIED HAND|JUVENILE ARTHRITIS, UNSPECIFIED, UNSPECIFIED HAND
C2901096|T046|M84.476A|ICD10CM|PATHOLOGICAL FRACTURE, UNSPECIFIED FOOT, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, UNSP FOOT, INIT ENCNTR FOR FRACTURE
C0153494|T191|C38.4|DMDICD10|MALIGNANT NEOPLASM OF PLEURA|BOESARTIGE NEUBILDUNG: PLEURA
C2890505|T037|T84.050A|ICD10CM|PERIPROSTHETIC OSTEOLYSIS OF INTERNAL PROSTHETIC RIGHT HIP JOINT, INITIAL ENCOUNTER|PERIPROSTH OSTEOLYSIS OF INTERNAL PROSTHETIC R HIP JT, INIT
C0153502|T191|C38.2|DMDICD10|MALIGNANT NEOPLASM OF POSTERIOR MEDIASTINUM|BOESARTIGE NEUBILDUNG: HINTERES MEDIASTINUM
C0153504|T191|C38.3|DMDICD10|MALIGNANT NEOPLASM OF MEDIASTINUM, PART UNSPECIFIED|BOESARTIGE NEUBILDUNG: MEDIASTINUM, TEIL NICHT NAEHER BEZEICHNET
C0346609|T191||ICD10CM|MALIGNANT NEOPLASM OF HEART
C0153501|T191|C38.1|DMDICD10|MALIGNANT NEOPLASM OF ANTERIOR MEDIASTINUM|BOESARTIGE NEUBILDUNG: VORDERES MEDIASTINUM
C0349042|T191|C38.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF HEART, MEDIASTINUM AND PLEURA|BOESARTIGE NEUBILDUNG: HERZ, MEDIASTINUM UND PLEURA, MEHRERE TEILBEREICHE UEBERLAPPEND
C2837993|T191|C43.39|ICD10CM|MALIGNANT MELANOMA OF OTHER PARTS OF FACE|MALIGNANT MELANOMA OF OTHER PARTS OF FACE
C2837991|T191|C43.30|ICD10CM|MALIGNANT MELANOMA OF UNSPECIFIED PART OF FACE|MALIGNANT MELANOMA OF UNSPECIFIED PART OF FACE
C2837992|T191|C43.31|ICD10CM|MALIGNANT MELANOMA OF NOSE|MALIGNANT MELANOMA OF NOSE
C4267937|T047|E08.3542|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, LEFT EYE|DIAB WITH PROLIF DIABETIC RTNOP WITH COMB DETACH, LEFT EYE
C4267938|T047|E08.3543|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, BILATERAL|DIABETES WITH PROLIF DIABETIC RTNOP WITH COMBINED DETACH, BI
C4267936|T047|E08.3541|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, RIGHT EYE|DIABETES WITH PROLIF DIABETIC RTNOP WITH COMB DETACH, R EYE
C2889905|T037|T82.318A|ICD10CM|BREAKDOWN (MECHANICAL) OF OTHER VASCULAR GRAFTS, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF OTHER VASCULAR GRAFTS, INIT ENCNTR
C4267939|T047|E08.3549|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH COMBINED TRACTION RETINAL DETACHMENT AND RHEGMATOGENOUS RETINAL DETACHMENT, UNSPECIFIED EYE|DIABETES WITH PROLIF DIABETIC RTNOP WITH COMB DETACH, UNSP
C2853782|T191|C81.98|ICD10CM|HODGKIN LYMPHOMA, UNSPECIFIED, LYMPH NODES OF MULTIPLE SITES|HODGKIN LYMPHOMA, UNSPECIFIED, LYMPH NODES OF MULTIPLE SITES
C2853783|T191|C81.99|ICD10CM|HODGKIN LYMPHOMA, UNSPECIFIED, EXTRANODAL AND SOLID ORGAN SITES|HODGKIN LYMPHOMA, UNSP, EXTRANODAL AND SOLID ORGAN SITES
C2853774|T191|C81.90|ICD10CM|HODGKIN LYMPHOMA, UNSPECIFIED, UNSPECIFIED SITE|HODGKIN LYMPHOMA, UNSPECIFIED, UNSPECIFIED SITE
C2853775|T191|C81.91|ICD10CM|HODGKIN LYMPHOMA, UNSPECIFIED, LYMPH NODES OF HEAD, FACE, AND NECK|HODGKIN LYMPHOMA, UNSP, LYMPH NODES OF HEAD, FACE, AND NECK
C2853776|T191|C81.92|ICD10CM|HODGKIN LYMPHOMA, UNSPECIFIED, INTRATHORACIC LYMPH NODES|HODGKIN LYMPHOMA, UNSPECIFIED, INTRATHORACIC LYMPH NODES
C2853777|T191|C81.93|ICD10CM|HODGKIN LYMPHOMA, UNSPECIFIED, INTRA-ABDOMINAL LYMPH NODES|HODGKIN LYMPHOMA, UNSPECIFIED, INTRA-ABDOMINAL LYMPH NODES
C2853778|T191|C81.94|ICD10CM|HODGKIN LYMPHOMA, UNSPECIFIED, LYMPH NODES OF AXILLA AND UPPER LIMB|HODGKIN LYMPHOMA, UNSP, LYMPH NODES OF AXILLA AND UPPER LIMB
C2853779|T191|C81.95|ICD10CM|HODGKIN LYMPHOMA, UNSPECIFIED, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|HODGKIN LYMPHOMA, UNSP, NODES OF ING REGION AND LOWER LIMB
C2853780|T191|C81.96|ICD10CM|HODGKIN LYMPHOMA, UNSPECIFIED, INTRAPELVIC LYMPH NODES|HODGKIN LYMPHOMA, UNSPECIFIED, INTRAPELVIC LYMPH NODES
C2853781|T191|C81.97|ICD10CM|HODGKIN LYMPHOMA, UNSPECIFIED, SPLEEN|HODGKIN LYMPHOMA, UNSPECIFIED, SPLEEN
C2977928|T191|C56.2|ICD10CM|MALIGNANT NEOPLASM OF LEFT OVARY|MALIGNANT NEOPLASM OF LEFT OVARY
C2842146|T191|C56.1|ICD10CM|MALIGNANT NEOPLASM OF RIGHT OVARY|MALIGNANT NEOPLASM OF RIGHT OVARY
C2842147|T191|C56.9|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED OVARY|MALIGNANT NEOPLASM OF UNSPECIFIED OVARY
C2885867|T037|T63.812A|ICD10CM|TOXIC EFFECT OF CONTACT WITH VENOMOUS FROG, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CONTACT W VENOMOUS FROG, SELF-HARM, INIT
C2832121|T037|S06.316S|ICD10CM|CONTUSION AND LACERATION OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|CONTUS/LAC R CEREB W LOC >24 HR W/O RET CONSC W SURV, SQLA
C2833480|T037|S12.44XB|ICD10CM|TYPE III TRAUMATIC SPONDYLOLISTHESIS OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE III TRAUM SPONDYLOLYSIS OF 5TH CERVCAL VERT, 7THB
C2977842|T037|S32.501B|ICD10CM|UNSPECIFIED FRACTURE OF RIGHT PUBIS, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF RIGHT PUBIS, INIT ENCNTR FOR OPEN FRACTURE
C2977841|T037|S32.501A|ICD10CM|UNSPECIFIED FRACTURE OF RIGHT PUBIS, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF RIGHT PUBIS, INIT FOR CLOS FX
C2832119|T037|S06.316A|ICD10CM|CONTUSION AND LACERATION OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|CONTUS/LAC R CEREB W LOC >24 HR W/O RET CONSC W SURV, INIT
C2885869|T037|T63.812S|ICD10CM|TOXIC EFFECT OF CONTACT WITH VENOMOUS FROG, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CONTACT W VENOMOUS FROG, SELF-HARM, SEQUELA
C2890471|T037|T84.038A|ICD10CM|MECHANICAL LOOSENING OF OTHER INTERNAL PROSTHETIC JOINT, INITIAL ENCOUNTER|MECHANICAL LOOSENING OF OTH INTERNAL PROSTHETIC JOINT, INIT
C2879440|T037|T46.2X2A|ICD10CM|POISONING BY OTHER ANTIDYSRHYTHMIC DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH ANTIDYSRHYTHMIC DRUGS, SELF-HARM, INIT
C2876594|T037|T36.2X2A|ICD10CM|POISONING BY CHLORAMPHENICOL GROUP, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY CHLORAMPHENICOL GROUP, SELF-HARM, INIT
C2834026|T037|S14.149D|ICD10CM|BROWN-SEQUARD SYNDROME AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|BROWN-SEQUARD SYND AT UNSP LEVEL OF CERV SPINAL CORD, SUBS
C0154222|T047|E31|DMDICD10|POLYGLANDULAR DYSFUNCTION, UNSPECIFIED|POLYGLANDULAERE DYSFUNKTION
C4268128|T047|E13.3219|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|OTH DIABETES WITH MILD NONP RTNOP WITH MACULAR EDEMA, UNSP
C2876596|T037|T36.2X2S|ICD10CM|POISONING BY CHLORAMPHENICOL GROUP, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY CHLORAMPHENICOL GROUP, SELF-HARM, SEQUELA
C4268126|T047|E13.3212|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|OTH DIAB WITH MILD NONP RTNOP WITH MACULAR EDEMA, LEFT EYE
C4268127|T047|E13.3213|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|OTH DIABETES WITH MILD NONP RTNOP WITH MACULAR EDEMA, BI
C0342556|T046|E31.1|DMDICD10|POLYGLANDULAR HYPERFUNCTION|POLYGLANDULAERE UEBERFUNKTION
C4268125|T047|E13.3211|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|OTH DIABETES WITH MILD NONP RTNOP WITH MACULAR EDEMA, R EYE
C2882365|T047|I63.312|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF LEFT MIDDLE CEREBRAL ARTERY|CEREBRAL INFRC DUE TO THOMBOS OF LEFT MIDDLE CEREBRAL ARTERY
C2882672|T047|I69.953|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING RIGHT NON-DOMINANT SIDE|HEMIPLGA FOL UNSP CEREBVASC DISEASE AFF RIGHT NONDOM SIDE
C2882364|T047|I63.311|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF RIGHT MIDDLE CEREBRAL ARTERY|CEREB INFRC DUE TO THOMBOS OF RIGHT MIDDLE CEREBRAL ARTERY
C2831994|T037|S06.1X5S|ICD10CM|TRAUMATIC CEREBRAL EDEMA WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, SEQUELA|TRAUM CEREBRAL EDEMA W LOC >24 HR W RET CONSC LEV, SEQUELA
C2882673|T047|I69.954|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING LEFT NON-DOMINANT SIDE|HEMIPLGA FOL UNSP CEREBVASC DISEASE AFF LEFT NONDOM SIDE
C2876134|T037|T31.31|ICD10CM|BURNS INVOLVING 30-39% OF BODY SURFACE WITH 10-19% THIRD DEGREE BURNS|BURNS OF 30-39% OF BODY SURFACE W 10-19% THIRD DEGREE BURNS
C0838553|T047|M46.91|ICD10CM|UNSPECIFIED INFLAMMATORY SPONDYLOPATHY, OCCIPITO-ATLANTO-AXIAL REGION|UNSP INFLAMMATORY SPONDYLOPATHY, OCCIPT-ATLAN-AX REGION
C0838561|T047|M46.90|ICD10CM|UNSPECIFIED INFLAMMATORY SPONDYLOPATHY, SITE UNSPECIFIED|UNSPECIFIED INFLAMMATORY SPONDYLOPATHY, SITE UNSPECIFIED
C0838555|T047|M46.93|ICD10CM|UNSPECIFIED INFLAMMATORY SPONDYLOPATHY, CERVICOTHORACIC REGION|UNSP INFLAMMATORY SPONDYLOPATHY, CERVICOTHORACIC REGION
C2882366|T047|I63.319|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF UNSPECIFIED MIDDLE CEREBRAL ARTERY|CEREBRAL INFRC DUE TO THOMBOS UNSP MIDDLE CEREBRAL ARTERY
C0838557|T047|M46.95|ICD10AM|UNSPECIFIED INFLAMMATORY SPONDYLOPATHY, THORACOLUMBAR REGION|UNSPECIFIED INFLAMMATORY SPONDYLOPATHY, THORACOLUMBAR REGION
C0838556|T047|M46.94|ICD10AM|UNSPECIFIED INFLAMMATORY SPONDYLOPATHY, THORACIC REGION|UNSPECIFIED INFLAMMATORY SPONDYLOPATHY, THORACIC REGION
C0838559|T047|M46.97|ICD10AM|UNSPECIFIED INFLAMMATORY SPONDYLOPATHY, LUMBOSACRAL REGION|UNSPECIFIED INFLAMMATORY SPONDYLOPATHY, LUMBOSACRAL REGION
C0838558|T047|M46.96|ICD10AM|UNSPECIFIED INFLAMMATORY SPONDYLOPATHY, LUMBAR REGION|UNSPECIFIED INFLAMMATORY SPONDYLOPATHY, LUMBAR REGION
C2873927|T047|E08.59|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH OTHER CIRCULATORY COMPLICATIONS|DIABETES DUE TO UNDERLYING CONDITION W OTH CIRCULATORY COMP
C2831992|T037|S06.1X5A|ICD10CM|TRAUMATIC CEREBRAL EDEMA WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, INITIAL ENCOUNTER|TRAUMATIC CEREBRAL EDEMA W LOC >24 HR W RET CONSC LEV, INIT
C2873926|T047|E08.52|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH DIABETIC PERIPHERAL ANGIOPATHY WITH GANGRENE|DIAB DUE TO UNDRL COND W DIABETIC PRPH ANGIOPATH W GANGRENE
C2873924|T047|E08.51|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH DIABETIC PERIPHERAL ANGIOPATHY WITHOUT GANGRENE|DIAB DUE TO UNDRL COND W DIAB PRPH ANGIOPATH W/O GANGRENE
C1409719|T047||ICD10CM|DISSEMINATED HERPESVIRAL DISEASE
C2833904|T037|S14.116S|ICD10CM|COMPLETE LESION AT C6 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|COMPLETE LESION AT C6 LEVEL OF CERVICAL SPINAL CORD, SEQUELA
C2857241|T037|S72.116C|ICD10CM|NONDISPLACED FRACTURE OF GREATER TROCHANTER OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF GREATER TROCHANTER OF UNSP FEMR, 7THC
C2857240|T037|S72.116B|ICD10CM|NONDISPLACED FRACTURE OF GREATER TROCHANTER OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF GREATER TROCHANTER OF UNSP FEMR, 7THB
C2857239|T037|S72.116A|ICD10CM|NONDISPLACED FRACTURE OF GREATER TROCHANTER OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF GREATER TROCHANTER OF UNSP FEMUR, INIT
C2833902|T037|S14.116A|ICD10CM|COMPLETE LESION AT C6 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION AT C6 LEVEL OF CERVICAL SPINAL CORD, INIT
C2833903|T037|S14.116D|ICD10CM|COMPLETE LESION AT C6 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION AT C6 LEVEL OF CERVICAL SPINAL CORD, SUBS
C4268294|T048|F19.27|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH PSYCHOACTIVE SUBSTANCE-INDUCED PERSISTING DEMENTIA|OTHER (OR UNKNOWN) SUBSTANCE USE DISORDER, SEVERE, WITH OTHER (OR UNKNOWN) SUBSTANCE INDUCED MAJOR NEUROCOGNITIVE DISORDER
C4268292|T048|F19.24|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH PSYCHOACTIVE SUBSTANCE-INDUCED MOOD DISORDER|OTHER (OR UNKNOWN) SUBSTANCE USE DISORDER, SEVERE, WITH OTHER (OR UNKNOWN) SUBSTANCE INDUCED DEPRESSIVE DISORDER
C2837503|T037|S32.018B|ICD10CM|OTHER FRACTURE OF FIRST LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF FIRST LUMBAR VERTEBRA, INIT FOR OPN FX
C2855855|T037|S68.022S|ICD10CM|PARTIAL TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF LEFT THUMB, SEQUELA|PARTIAL TRAUMATIC MCP AMPUTATION OF LEFT THUMB, SEQUELA
C2889969|T037|T82.398A|ICD10CM|OTHER MECHANICAL COMPLICATION OF OTHER VASCULAR GRAFTS, INITIAL ENCOUNTER|MECH COMPL OF OTHER VASCULAR GRAFTS, INITIAL ENCOUNTER
C2889644|T047|M08.959|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, UNSPECIFIED HIP|JUVENILE ARTHRITIS, UNSPECIFIED, UNSPECIFIED HIP
C2860025|T037|S78.911S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT HIP AND THIGH, LEVEL UNSPECIFIED, SEQUELA|COMPLETE TRAUM AMP OF R HIP AND THIGH, LEVEL UNSP, SEQUELA
C2859986|T037|S78.021S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT RIGHT HIP JOINT, SEQUELA|PARTIAL TRAUMATIC AMPUTATION AT RIGHT HIP JOINT, SEQUELA
C2889643|T047|M08.952|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, LEFT HIP|JUVENILE ARTHRITIS, UNSPECIFIED, LEFT HIP
C2889642|T047|M08.951|ICD10CM|JUVENILE ARTHRITIS, UNSPECIFIED, RIGHT HIP|JUVENILE ARTHRITIS, UNSPECIFIED, RIGHT HIP
C2859985|T037|S78.021D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT RIGHT HIP JOINT, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION AT RIGHT HIP JOINT, SUBS ENCNTR
C2901823|T047|M86.222|ICD10CM|SUBACUTE OSTEOMYELITIS, LEFT HUMERUS|SUBACUTE OSTEOMYELITIS, LEFT HUMERUS
C2901822|T047|M86.221|ICD10CM|SUBACUTE OSTEOMYELITIS, RIGHT HUMERUS|SUBACUTE OSTEOMYELITIS, RIGHT HUMERUS
C2879570|T037|T46.7X2S|ICD10CM|POISONING BY PERIPHERAL VASODILATORS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY PERIPHERAL VASODILATORS, SELF-HARM, SEQUELA
C2884018|T037|T51.2X2A|ICD10CM|TOXIC EFFECT OF 2-PROPANOL, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF 2-PROPANOL, INTENTIONAL SELF-HARM, INIT
C2890418|T037|T84.018A|ICD10CM|BROKEN INTERNAL JOINT PROSTHESIS, OTHER SITE, INITIAL ENCOUNTER|BROKEN INTERNAL JOINT PROSTHESIS, OTHER SITE, INIT ENCNTR
C2901824|T047|M86.229|ICD10CM|SUBACUTE OSTEOMYELITIS, UNSPECIFIED HUMERUS|SUBACUTE OSTEOMYELITIS, UNSPECIFIED HUMERUS
C2853901|T191|C83.18|ICD10CM|MANTLE CELL LYMPHOMA, LYMPH NODES OF MULTIPLE SITES|MANTLE CELL LYMPHOMA, LYMPH NODES OF MULTIPLE SITES
C0348826|T047|D86.2|DMDICD10|SARCOIDOSIS OF LUNG WITH SARCOIDOSIS OF LYMPH NODES|SARKOIDOSE DER LUNGE MIT SARKOIDOSE DER LYMPHKNOTEN
C0036205|T047|D86.0|DMDICD10|SARCOIDOSIS OF LUNG|SARKOIDOSE DER LUNGE
C2855989|T037|S68.521S|ICD10CM|PARTIAL TRAUMATIC TRANSPHALANGEAL AMPUTATION OF RIGHT THUMB, SEQUELA|PARTIAL TRAUMATIC TRNSPHAL AMPUTATION OF R THM, SEQUELA
C2835355|T037|S22.058A|ICD10CM|OTHER FRACTURE OF T5-T6 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF T5-T6 VERTEBRA, INIT FOR CLOS FX
C2835356|T037|S22.058B|ICD10CM|OTHER FRACTURE OF T5-T6 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF T5-T6 VERTEBRA, INIT FOR OPN FX
C0151517|T047|I44.2|DMDICD10|ATRIOVENTRICULAR BLOCK, COMPLETE|ATRIOVENTRIKULAERER BLOCK 3. GRADES
C2890032|T037|T82.520A|ICD10CM|DISPLACEMENT OF SURGICALLY CREATED ARTERIOVENOUS FISTULA, INITIAL ENCOUNTER|DISPLACEMENT OF SURGICALLY CREATED AV FISTULA, INIT
C0270942|T047||ICD10CM|MYASTHENIA GRAVIS WITH (ACUTE) EXACERBATION
C1260409|T047||ICD10CM|MYASTHENIA GRAVIS WITHOUT (ACUTE) EXACERBATION
C2901459|T046|M84.642A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, LEFT HAND, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, LEFT HAND, INIT FOR FX
C2835802|T037|S24.132D|ICD10CM|ANTERIOR CORD SYNDROME AT T2-T6 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|ANTERIOR CORD SYNDROME AT T2-T6, SUBS
C2890003|T037|T82.511A|ICD10CM|BREAKDOWN (MECHANICAL) OF SURGICALLY CREATED ARTERIOVENOUS SHUNT, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF SURGICALLY CREATED AV SHUNT, INIT
C2835835|T037|S24.149D|ICD10CM|BROWN-SEQUARD SYNDROME AT UNSPECIFIED LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|BROWN-SEQUARD SYND AT UNSP LEVEL OF THOR SPINAL CORD, SUBS
C4270292|T046|T83.411A|ICD10CM|BREAKDOWN (MECHANICAL) OF IMPLANTED TESTICULAR PROSTHESIS, INITIAL ENCOUNTER|BREAKDOWN OF IMPLANTED TESTICULAR PROSTHESIS, INIT
C2835801|T037|S24.132A|ICD10CM|ANTERIOR CORD SYNDROME AT T2-T6 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|ANTERIOR CORD SYNDROME AT T2-T6, INIT
C2835834|T037|S24.149A|ICD10CM|BROWN-SEQUARD SYNDROME AT UNSPECIFIED LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|BROWN-SEQUARD SYND AT UNSP LEVEL OF THOR SPINAL CORD, INIT
C2835836|T037|S24.149S|ICD10CM|BROWN-SEQUARD SYNDROME AT UNSPECIFIED LEVEL OF THORACIC SPINAL CORD, SEQUELA|BROWN-SEQUARD SYND AT UNSP LEVEL OF THOR SPINAL CORD, SQLA
C2835803|T037|S24.132S|ICD10CM|ANTERIOR CORD SYNDROME AT T2-T6 LEVEL OF THORACIC SPINAL CORD, SEQUELA|ANTERIOR CORD SYNDROME AT T2-T6, SEQUELA
C2833953|T037|S14.129S|ICD10CM|CENTRAL CORD SYNDROME AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, SEQUELA|CENTRAL CORD SYND AT UNSP LEVEL OF CERV SPINAL CORD, SEQUELA
C2884203|T037|T53.0X2S|ICD10CM|TOXIC EFFECT OF CARBON TETRACHLORIDE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CARBON TETRACHLORIDE, SELF-HARM, SEQUELA
C2879128|T037|T45.4X2S|ICD10CM|POISONING BY IRON AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY IRON AND ITS COMPOUNDS, SELF-HARM, SEQUELA
C2884201|T037|T53.0X2A|ICD10CM|TOXIC EFFECT OF CARBON TETRACHLORIDE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CARBON TETRACHLORIDE, SELF-HARM, INIT
C2833532|T037|S12.530A|ICD10CM|UNSPECIFIED TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP TRAUM DISPL SPONDYLOLYSIS OF SIXTH CERVCAL VERT, INIT
C2879126|T037|T45.4X2A|ICD10CM|POISONING BY IRON AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY IRON AND ITS COMPOUNDS, SELF-HARM, INIT
C2833533|T037|S12.530B|ICD10CM|UNSPECIFIED TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP TRAUM DISPL SPONDYLOLYSIS OF SIXTH CERVCAL VERT, 7THB
C2869776|T037|S98.029A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED FOOT AT ANKLE LEVEL, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP OF UNSP FOOT AT ANKLE LEVEL, INIT
C2833884|T037|S14.111S|ICD10CM|COMPLETE LESION AT C1 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|COMPLETE LESION AT C1 LEVEL OF CERVICAL SPINAL CORD, SEQUELA
C2833472|T037|S12.431A|ICD10CM|UNSPECIFIED TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP TRAUM NONDISP SPONDYLOLYSIS OF FIFTH CERVCAL VERT, INIT
C2833473|T037|S12.431B|ICD10CM|UNSPECIFIED TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP TRAUM NONDISP SPONDYLOLYSIS OF 5TH CERVCAL VERT, 7THB
C2901941|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF LEFT HUMERUS
C2889163|T047|M05.179|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT|RHEU LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP ANK/FT
C2882729|T047|I70.248|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF LEFT LEG WITH ULCERATION OF OTHER PART OF LOWER LEFT LEG|ATHSCL NATIVE ART OF LEFT LEG W ULCER OTH PRT LOWER LEFT LEG
C2882730|T047|I70.249|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF LEFT LEG WITH ULCERATION OF UNSPECIFIED SITE|ATHSCL NATIVE ARTERIES OF LEFT LEG W ULCERATION OF UNSP SITE
C2845879|T191|C62.91|ICD10CM|MALIGNANT NEOPLASM OF RIGHT TESTIS, UNSPECIFIED WHETHER DESCENDED OR UNDESCENDED|MALIG NEOPLM OF RIGHT TESTIS, UNSP DESCENDED OR UNDESCENDED
C2845878|T191|C62.90|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED TESTIS, UNSPECIFIED WHETHER DESCENDED OR UNDESCENDED|MALIG NEOPLASM OF UNSP TESTIS, UNSP DESCENDED OR UNDESCENDED
C2845880|T191|C62.92|ICD10CM|MALIGNANT NEOPLASM OF LEFT TESTIS, UNSPECIFIED WHETHER DESCENDED OR UNDESCENDED|MALIG NEOPLASM OF LEFT TESTIS, UNSP DESCENDED OR UNDESCENDED
C2882722|T047|I70.241|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF LEFT LEG WITH ULCERATION OF THIGH|ATHSCL NATIVE ARTERIES OF LEFT LEG W ULCERATION OF THIGH
C2882723|T047|I70.242|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF LEFT LEG WITH ULCERATION OF CALF|ATHSCL NATIVE ARTERIES OF LEFT LEG W ULCERATION OF CALF
C2882724|T047|I70.243|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF LEFT LEG WITH ULCERATION OF ANKLE|ATHSCL NATIVE ARTERIES OF LEFT LEG W ULCERATION OF ANKLE
C2901999|T046|M87.137|ICD10CM|OSTEONECROSIS DUE TO DRUGS OF RIGHT CARPUS|OSTEONECROSIS DUE TO DRUGS OF RIGHT CARPUS
C2891230|T037|T85.79XA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO OTHER INTERNAL PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO OTH INT PROSTH DEV/GRFT, INIT
C2884742|T037|T58.02XA|ICD10CM|TOXIC EFFECT OF CARBON MONOXIDE FROM MOTOR VEHICLE EXHAUST, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFF OF CARB MONX FROM MTR VEH EXHAUST, SLF-HRM, INIT
C2878484|T037|T43.4X2S|ICD10CM|POISONING BY BUTYROPHENONE AND THIOTHIXENE NEUROLEPTICS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY BUTYROPHEN/THIOTHIXEN NEUROLEPTC, SLF-HRM, SEQUELA
C4268631|T047|K55.059|ICD10CM|ACUTE (REVERSIBLE) ISCHEMIA OF INTESTINE, PART AND EXTENT UNSPECIFIED|ACUTE ISCHEMIA OF INTESTINE, PART AND EXTENT UNSPECIFIED
C3264203|T047|H40.1232|ICD10CM|LOW-TENSION GLAUCOMA, BILATERAL, MODERATE STAGE|LOW-TENSION GLAUCOMA, BILATERAL, MODERATE STAGE
C4268630|T047|K55.052|ICD10CM|DIFFUSE ACUTE (REVERSIBLE) ISCHEMIA OF INTESTINE, PART UNSPECIFIED|DIFFUSE ACUTE ISCHEMIA OF INTESTINE, PART UNSPECIFIED
C4268629|T047|K55.051|ICD10CM|FOCAL (SEGMENTAL) ACUTE (REVERSIBLE) ISCHEMIA OF INTESTINE, PART UNSPECIFIED|FOCAL ACUTE ISCHEMIA OF INTESTINE, PART UNSPECIFIED
C2885322|T037|T63.012A|ICD10CM|TOXIC EFFECT OF RATTLESNAKE VENOM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF RATTLESNAKE VENOM, SELF-HARM, INIT
C2858149|T037|S72.362B|ICD10CM|DISPLACED SEGMENTAL FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL SEG FX SHAFT OF L FEMUR, INIT FOR OPN FX TYPE I/2
C2858150|T037|S72.362C|ICD10CM|DISPLACED SEGMENTAL FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL SEG FX SHAFT OF L FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2858148|T037|S72.362A|ICD10CM|DISPLACED SEGMENTAL FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED SEGMENTAL FRACTURE OF SHAFT OF LEFT FEMUR, INIT
C2874939|T048|F40.228|ICD10CM|OTHER NATURAL ENVIRONMENT TYPE PHOBIA|OTHER NATURAL ENVIRONMENT TYPE PHOBIA
C2869777|T037|S98.029D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED FOOT AT ANKLE LEVEL, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMP OF UNSP FOOT AT ANKLE LEVEL, SUBS
C0558207|T048||ICD10CM|FEAR OF THUNDERSTORMS
C2885324|T037|T63.012S|ICD10CM|TOXIC EFFECT OF RATTLESNAKE VENOM, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF RATTLESNAKE VENOM, SELF-HARM, SEQUELA
C2877741|T037|T40.692S|ICD10CM|POISONING BY OTHER NARCOTICS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTHER NARCOTICS, INTENTIONAL SELF-HARM, SEQUELA
C3264181|T047|H40.10X0|ICD10CM|UNSPECIFIED OPEN-ANGLE GLAUCOMA, STAGE UNSPECIFIED|UNSPECIFIED OPEN-ANGLE GLAUCOMA, STAGE UNSPECIFIED
C3264182|T047|H40.10X1|ICD10CM|UNSPECIFIED OPEN-ANGLE GLAUCOMA, MILD STAGE|UNSPECIFIED OPEN-ANGLE GLAUCOMA, MILD STAGE
C3264183|T047|H40.10X2|ICD10CM|UNSPECIFIED OPEN-ANGLE GLAUCOMA, MODERATE STAGE|UNSPECIFIED OPEN-ANGLE GLAUCOMA, MODERATE STAGE
C3264184|T047|H40.10X3|ICD10CM|UNSPECIFIED OPEN-ANGLE GLAUCOMA, SEVERE STAGE|UNSPECIFIED OPEN-ANGLE GLAUCOMA, SEVERE STAGE
C3264185|T047|H40.10X4|ICD10CM|UNSPECIFIED OPEN-ANGLE GLAUCOMA, INDETERMINATE STAGE|UNSPECIFIED OPEN-ANGLE GLAUCOMA, INDETERMINATE STAGE
C2869804|T037|S98.129S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED GREAT TOE, SEQUELA|PARTIAL TRAUMATIC AMPUTATION OF UNSP GREAT TOE, SEQUELA
C2521695|T060|C715|ICD10PCS|MALIGNANT NEOPLASM OF CEREBRAL VENTRICLE|NUCLEAR MEDICINE @ LYMPHATIC AND HEMATOLOGIC SYSTEM @ PLANAR NUCLEAR MEDICINE IMAGING @ LYMPHATICS, HEAD AND NECK
C0153638|T191|C71.4|DMDICD10|MALIGNANT NEOPLASM OF OCCIPITAL LOBE|BOESARTIGE NEUBILDUNG: OKZIPITALLAPPEN
C2845928|T191|C71.7|ICD10CM|MALIGNANT NEOPLASM OF BRAIN STEM|MALIGNANT NEOPLASM OF FOURTH CEREBRAL VENTRICLE
C0153640|T191|C71.6|DMDICD10|MALIGNANT NEOPLASM OF CEREBELLUM|BOESARTIGE NEUBILDUNG: ZEREBELLUM
C0153635|T191|C71.1|DMDICD10|MALIGNANT NEOPLASM OF FRONTAL LOBE|BOESARTIGE NEUBILDUNG: FRONTALLAPPEN
C2521683|T060|C710|ICD10PCS|MALIGNANT NEOPLASM OF CEREBRUM, EXCEPT LOBES AND VENTRICLES|NUCLEAR MEDICINE @ LYMPHATIC AND HEMATOLOGIC SYSTEM @ PLANAR NUCLEAR MEDICINE IMAGING @ BONE MARROW
C2521735|T060|C713|ICD10PCS|MALIGNANT NEOPLASM OF PARIETAL LOBE|NUCLEAR MEDICINE @ LYMPHATIC AND HEMATOLOGIC SYSTEM @ PLANAR NUCLEAR MEDICINE IMAGING @ BLOOD
C2521690|T060|C712|ICD10PCS|MALIGNANT NEOPLASM OF TEMPORAL LOBE|NUCLEAR MEDICINE @ LYMPHATIC AND HEMATOLOGIC SYSTEM @ PLANAR NUCLEAR MEDICINE IMAGING @ SPLEEN
C0153633|T191|C71.9|DMDICD10|MALIGNANT NEOPLASM OF BRAIN, UNSPECIFIED|BOESARTIGE NEUBILDUNG: GEHIRN, NICHT NAEHER BEZEICHNET
C0496837|T191|C71.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF BRAIN|BOESARTIGE NEUBILDUNG: GEHIRN, MEHRERE TEILBEREICHE UEBERLAPPEND
C2888666|T047|L97.213|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT CALF WITH NECROSIS OF MUSCLE|NON-PRS CHRONIC ULCER OF RIGHT CALF W NECROSIS OF MUSCLE
C2888665|T047|L97.212|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT CALF WITH FAT LAYER EXPOSED|NON-PRESSURE CHRONIC ULCER OF RIGHT CALF W FAT LAYER EXPOSED
C2888664|T047|L97.211|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT CALF LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHRONIC ULCER OF RIGHT CALF LIMITED TO BRKDWN SKIN
C2885951|T037|T64.02XS|ICD10CM|TOXIC EFFECT OF AFLATOXIN, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF AFLATOXIN, INTENTIONAL SELF-HARM, SEQUELA
C4509288|T047|L97.216|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT CALF WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULCER OF R CALF WITH BONE INVL W/O EVD OF NECR
C4509287|T047|L97.215|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT CALF WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULCER OF R CALF WITH MSL INVL W/O EVD OF NECR
C2888667|T047|L97.214|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT CALF WITH NECROSIS OF BONE|NON-PRESSURE CHRONIC ULCER OF RIGHT CALF W NECROSIS OF BONE
C2835788|T037|S24.114A|ICD10CM|COMPLETE LESION AT T11-T12 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|COMPLETE LESION AT T11-T12, INIT
C2888668|T047|L97.219|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT CALF WITH UNSPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF RIGHT CALF WITH UNSP SEVERITY
C4509289|T047|L97.218|ICD10CM|NON-PRESSURE CHRONIC ULCER OF RIGHT CALF WITH OTHER SPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OF RIGHT CALF WITH OTH SEVERITY
C2835789|T037|S24.114D|ICD10CM|COMPLETE LESION AT T11-T12 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION AT T11-T12, SUBS
C2857977|T037|S72.344B|ICD10CM|NONDISPLACED SPIRAL FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP SPIRAL FX SHAFT OF R FEMUR, INIT FOR OPN FX TYPE I/2
C2857978|T037|S72.344C|ICD10CM|NONDISPLACED SPIRAL FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP SPIRAL FX SHAFT OF R FEMR, 7THC
C2885949|T037|T64.02XA|ICD10CM|TOXIC EFFECT OF AFLATOXIN, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF AFLATOXIN, INTENTIONAL SELF-HARM, INIT
C2857976|T037|S72.344A|ICD10CM|NONDISPLACED SPIRAL FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED SPIRAL FRACTURE OF SHAFT OF RIGHT FEMUR, INIT
C2877384|T037|T39.1X2S|ICD10CM|POISONING BY 4-AMINOPHENOL DERIVATIVES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY 4-AMINOPHENOL DERIVATIVES, SELF-HARM, SEQUELA
C2835790|T037|S24.114S|ICD10CM|COMPLETE LESION AT T11-T12 LEVEL OF THORACIC SPINAL CORD, SEQUELA|COMPLETE LESION AT T11-T12, SEQUELA
C2838416|T037|S32.602B|ICD10CM|UNSPECIFIED FRACTURE OF LEFT ISCHIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF LEFT ISCHIUM, INIT ENCNTR FOR OPEN FRACTURE
C2838415|T037|S32.602A|ICD10CM|UNSPECIFIED FRACTURE OF LEFT ISCHIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF LEFT ISCHIUM, INIT FOR CLOS FX
C2876718|T037|T36.7X2A|ICD10CM|POISONING BY ANTIFUNGAL ANTIBIOTICS, SYSTEMICALLY USED, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ANTIFUNGAL ANTIBIOT, SYS USED, SELF-HARM, INIT
C2837957|T191|C34.80|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF UNSPECIFIED BRONCHUS AND LUNG|MALIGNANT NEOPLASM OF OVRLP SITES OF UNSP BRONCHUS AND LUNG
C2838194|T037|S32.453B|ICD10CM|DISPLACED TRANSVERSE FRACTURE OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISPLACED TRANSVERSE FX UNSP ACETABULUM, INIT FOR OPN FX
C2838193|T037|S32.453A|ICD10CM|DISPLACED TRANSVERSE FRACTURE OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED TRANSVERSE FRACTURE OF UNSP ACETABULUM, INIT
C2890608|T037|T84.117A|ICD10CM|BREAKDOWN (MECHANICAL) OF INTERNAL FIXATION DEVICE OF BONE OF LEFT LOWER LEG, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF INT FIX OF BONE OF L LOW LEG, INIT
C2889062|T047|M02.341|ICD10CM|REITER'S DISEASE, RIGHT HAND|REITER'S DISEASE, RIGHT HAND
C2889063|T047|M02.342|ICD10CM|REITER'S DISEASE, LEFT HAND|REITER'S DISEASE, LEFT HAND
C2889064|T047|M02.349|ICD10CM|REITER'S DISEASE, UNSPECIFIED HAND|REITER'S DISEASE, UNSPECIFIED HAND
C2869802|T037|S98.129A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED GREAT TOE, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF UNSP GREAT TOE, INIT ENCNTR
C0477596|T047|M36.8|DMDICD10|SYSTEMIC DISORDERS OF CONNECTIVE TISSUE IN OTHER DISEASES CLASSIFIED ELSEWHERE|SYSTEMKRANKHEITEN DES BINDEGEWEBES BEI SONSTIGEN ANDERENORTS KLASSIFIZIERTEN KRANKHEITEN
C2853840|T191|C82.52|ICD10CM|DIFFUSE FOLLICLE CENTER LYMPHOMA, INTRATHORACIC LYMPH NODES|DIFFUSE FOLLICLE CENTER LYMPHOMA, INTRATHORACIC LYMPH NODES
C3264037|T047|G43.A0|ICD10CM|CYCLICAL VOMITING, NOT INTRACTABLE|CYCLICAL VOMITING, WITHOUT REFRACTORY MIGRAINE
C3264038|T047|G43.A1|ICD10CM|CYCLICAL VOMITING, INTRACTABLE|CYCLICAL VOMITING, WITH REFRACTORY MIGRAINE
C0409990|T047|M36.0|DMDICD10|DERMATO(POLY)MYOSITIS IN NEOPLASTIC DISEASE|DERMATOMYOSITIS-POLYMYOSITIS BEI NEUBILDUNGEN
C3648005|T191|C82.51|ICD10CM|DIFFUSE FOLLICLE CENTER LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK|DIFFUSE FOLICL CENTER LYMPH, NODES OF HEAD, FACE, AND NECK
C2845956|T191|C76.52|ICD10CM|MALIGNANT NEOPLASM OF LEFT LOWER LIMB|MALIGNANT NEOPLASM OF LEFT LOWER LIMB
C2845954|T191|C76.50|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED LOWER LIMB|MALIGNANT NEOPLASM OF UNSPECIFIED LOWER LIMB
C2845955|T191|C76.51|ICD10CM|MALIGNANT NEOPLASM OF RIGHT LOWER LIMB|MALIGNANT NEOPLASM OF RIGHT LOWER LIMB
C2877228|T037|T38.812S|ICD10CM|POISONING BY ANTERIOR PITUITARY [ADENOHYPOPHYSEAL] HORMONES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ANTERIOR PITUITARY HORMONES, SELF-HARM, SEQUELA
C2858784|T037|S72.453C|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL SUPRCNDL FX W/O INTRCNDL EXTN LOW END UNSP FEMR, 7THC
C2858783|T037|S72.453B|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL SUPRCNDL FX W/O INTRCNDL EXTN LOW END UNSP FEMR, 7THB
C2858782|T037|S72.453A|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPL SUPRCNDL FX W/O INTRCNDL EXTN LOW END UNSP FEMR, INIT
C2877226|T037|T38.812A|ICD10CM|POISONING BY ANTERIOR PITUITARY [ADENOHYPOPHYSEAL] HORMONES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ANTERIOR PITUITARY HORMONES, SELF-HARM, INIT
C2886052|T037|T65.292S|ICD10CM|TOXIC EFFECT OF OTHER TOBACCO AND NICOTINE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF TOBACCO AND NICOTINE, SELF-HARM, SEQUELA
C2874218|T047|E44.0|ICD10CM|MODERATE PROTEIN-CALORIE MALNUTRITION|MODERATE PROTEIN-CALORIE MALNUTRITION
C2891286|T037|T86.819|ICD10CM|UNSPECIFIED COMPLICATION OF LUNG TRANSPLANT|UNSPECIFIED COMPLICATION OF LUNG TRANSPLANT
C2891285|T037|T86.818|ICD10CM|OTHER COMPLICATIONS OF LUNG TRANSPLANT|OTHER COMPLICATIONS OF LUNG TRANSPLANT
C2877407|T037|T39.2X2A|ICD10CM|POISONING BY PYRAZOLONE DERIVATIVES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY PYRAZOLONE DERIVATIVES, SELF-HARM, INIT
C2891284|T046||ICD10CM|LUNG TRANSPLANT INFECTION
C1404116|T046||ICD10CM|LUNG TRANSPLANT FAILURE
C0729958|T046|T86.810|ICD10CM|LUNG TRANSPLANT REJECTION|LUNG TRANSPLANT REJECTION
C2886050|T037|T65.292A|ICD10CM|TOXIC EFFECT OF OTHER TOBACCO AND NICOTINE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF TOBACCO AND NICOTINE, SELF-HARM, INIT
C3264046|T047|G71.0|ICD10CM|MUSCULAR DYSTROPHY|CONGENITAL MUSCULAR DYSTROPHY WITH SPECIFIC MORPHOLOGICAL ABNORMALITIES OF THE MUSCLE FIBER
C0869052|T047|G71.3|DMDICD10|MITOCHONDRIAL MYOPATHY, NOT ELSEWHERE CLASSIFIED|MITOCHONDRIALE MYOPATHIE, ANDERENORTS NICHT KLASSIFIZIERT
C2875316|T019|G71.2|ICD10CM|CONGENITAL MYOPATHIES|MYOTUBULAR (CENTRONUCLEAR) MYOPATHY
C2875076|T047|G40.001|ICD10CM|LOCALIZATION-RELATED (FOCAL) (PARTIAL) IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SEIZURES OF LOCALIZED ONSET, NOT INTRACTABLE, WITH STATUS EPILEPTICUS|LOCAL-REL IDIO EPI W SEIZ OF LOC ONST, NOT NTRCT, W STAT EPI
C2833824|T047|B97.35|ICD10CM|HUMAN IMMUNODEFICIENCY VIRUS, TYPE 2 [HIV 2] AS THE CAUSE OF DISEASES CLASSIFIED ELSEWHERE|HIV 2 AS THE CAUSE OF DISEASES CLASSIFIED ELSEWHERE
C1399469|T047||ICD10CM|PRIMARY DISORDER OF MUSCLE, UNSPECIFIED
C2874798|T048|F19.150|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE ABUSE WITH PSYCHOACTIVE SUBSTANCE-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|OTH PSYCHOACTV SUBSTANCE ABUSE W PSYCH DISORDER W DELUSIONS
C2875077|T047|G40.009|ICD10CM|LOCALIZATION-RELATED (FOCAL) (PARTIAL) IDIOPATHIC EPILEPSY AND EPILEPTIC SYNDROMES WITH SEIZURES OF LOCALIZED ONSET, NOT INTRACTABLE, WITHOUT STATUS EPILEPTICUS|LOCAL-REL IDIO EPI W SEIZ OF LOC ONST,NOT NTRCT,W/O STAT EPI
C2874799|T048|F19.151|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE ABUSE WITH PSYCHOACTIVE SUBSTANCE-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|OTH PSYCHOACTV SUBSTANCE ABUSE W PSYCH DISORDER W HALLUCIN
C4509308|T047|L97.425|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT HEEL AND MIDFOOT WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OF L HEEL/MIDFT W MSL INVL W/O EVD OF NECR
C2835169|T037|S22.002B|ICD10CM|UNSTABLE BURST FRACTURE OF UNSPECIFIED THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSTABLE BURST FX UNSP THOR VERTEBRA, INIT FOR OPN FX
C2890571|T037|T84.098A|ICD10CM|OTHER MECHANICAL COMPLICATION OF OTHER INTERNAL JOINT PROSTHESIS, INITIAL ENCOUNTER|MECH COMPL OF OTHER INTERNAL JOINT PROSTHESIS, INIT ENCNTR
C2888709|T047|L97.421|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT HEEL AND MIDFOOT LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHR ULCER OF LEFT HEEL AND MIDFT LMT TO BRKDWN SKIN
C2901386|T046|M84.619A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, UNSPECIFIED SHOULDER, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, UNSP SHOULDER, INIT
C2888711|T047|L97.423|ICD10CM|NON-PRESSURE CHRONIC ULCER OF LEFT HEEL AND MIDFOOT WITH NECROSIS OF MUSCLE|NON-PRS CHR ULCER OF LEFT HEEL AND MIDFOOT W NECROS MUSCLE
C4268169|T047|E13.3551|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, RIGHT EYE|OTH DIABETES WITH STABLE PROLIF DIABETIC RTNOP, RIGHT EYE
C2905791|T037|X82.0XXD|ICD10CM|INTENTIONAL COLLISION OF MOTOR VEHICLE WITH OTHER MOTOR VEHICLE, SUBSEQUENT ENCOUNTER|INTENTIONAL COLLISION OF MOTOR VEHICLE W MTR VEH, SUBS
C4268171|T047|E13.3553|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, BILATERAL|OTH DIABETES WITH STABLE PROLIF DIABETIC RTNOP, BILATERAL
C4268170|T047|E13.3552|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, LEFT EYE|OTH DIABETES WITH STABLE PROLIF DIABETIC RTNOP, LEFT EYE
C2905790|T037|X82.0XXA|ICD10CM|INTENTIONAL COLLISION OF MOTOR VEHICLE WITH OTHER MOTOR VEHICLE, INITIAL ENCOUNTER|INTENTIONAL COLLISION OF MOTOR VEHICLE W MTR VEH, INIT
C4268172|T047|E13.3559|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH STABLE PROLIFERATIVE DIABETIC RETINOPATHY, UNSPECIFIED EYE|OTH DIABETES WITH STABLE PROLIF DIABETIC RETINOPATHY, UNSP
C2890875|T037|T84.624A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL FIXATION DEVICE OF RIGHT FIBULA, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INT FIX OF RIGHT FIBULA, INIT
C0838510|T047|M46.28|ICD10AM|OSTEOMYELITIS OF VERTEBRA, SACRAL AND SACROCOCCYGEAL REGION|OSTEOMYELITIS OF VERTEBRA, SACRAL AND SACROCOCCYGEAL REGION
C2905792|T037|X82.0XXS|ICD10CM|INTENTIONAL COLLISION OF MOTOR VEHICLE WITH OTHER MOTOR VEHICLE, SEQUELA|INTENTIONAL COLLISION OF MOTOR VEHICLE W MTR VEH, SEQUELA
C2889205|T047|M05.322|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT ELBOW|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF L ELBOW
C2853944|T191|C83.89|ICD10CM|OTHER NON-FOLLICULAR LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES|OTH NON-FOLLIC LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES
C2853943|T191|C83.88|ICD10CM|OTHER NON-FOLLICULAR LYMPHOMA, LYMPH NODES OF MULTIPLE SITES|OTHER NON-FOLLICULAR LYMPHOMA, LYMPH NODES OF MULTIPLE SITES
C2893649|T047|M12.062|ICD10CM|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], LEFT KNEE|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], LEFT KNEE
C2853940|T191|C83.85|ICD10CM|OTHER NON-FOLLICULAR LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|OTH NON-FOLLIC LYMPHOMA, NODES OF ING REGION AND LOWER LIMB
C2853939|T191|C83.84|ICD10CM|OTHER NON-FOLLICULAR LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB|OTH NON-FOLLIC LYMPHOMA, NODES OF AXILLA AND UPPER LIMB
C2853942|T191|C83.87|ICD10CM|OTHER NON-FOLLICULAR LYMPHOMA, SPLEEN|OTHER NON-FOLLICULAR LYMPHOMA, SPLEEN
C2853941|T191|C83.86|ICD10CM|OTHER NON-FOLLICULAR LYMPHOMA, INTRAPELVIC LYMPH NODES|OTHER NON-FOLLICULAR LYMPHOMA, INTRAPELVIC LYMPH NODES
C2853936|T191|C83.81|ICD10CM|OTHER NON-FOLLICULAR LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK|OTH NON-FOLLIC LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK
C2853935|T191|C83.80|ICD10CM|OTHER NON-FOLLICULAR LYMPHOMA, UNSPECIFIED SITE|OTHER NON-FOLLICULAR LYMPHOMA, UNSPECIFIED SITE
C2853938|T191|C83.83|ICD10CM|OTHER NON-FOLLICULAR LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES|OTHER NON-FOLLICULAR LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES
C2853937|T191|C83.82|ICD10CM|OTHER NON-FOLLICULAR LYMPHOMA, INTRATHORACIC LYMPH NODES|OTHER NON-FOLLICULAR LYMPHOMA, INTRATHORACIC LYMPH NODES
C2832596|T037|S06.821S|ICD10CM|INJURY OF LEFT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|INJ L INT CRTD, INTCR W LOC OF 30 MINUTES OR LESS, SEQUELA
C2891187|T037|T85.631S|ICD10CM|LEAKAGE OF INTRAPERITONEAL DIALYSIS CATHETER, SEQUELA|LEAKAGE OF INTRAPERITONEAL DIALYSIS CATHETER, SEQUELA
C2885175|T037|T61.782S|ICD10CM|OTHER SHELLFISH POISONING, INTENTIONAL SELF-HARM, SEQUELA|OTHER SHELLFISH POISONING, INTENTIONAL SELF-HARM, SEQUELA
C0837061|T047|E13.11|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH KETOACIDOSIS WITH COMA|OTH DIABETES MELLITUS WITH KETOACIDOSIS WITH COMA
C0837060|T047|E13.10|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH KETOACIDOSIS WITHOUT COMA|OTH DIABETES MELLITUS WITH KETOACIDOSIS WITHOUT COMA
C2854083|T191|C90.30|ICD10CM|SOLITARY PLASMACYTOMA NOT HAVING ACHIEVED REMISSION|SOLITARY PLASMACYTOMA NOT HAVING ACHIEVED REMISSION
C2854084|T191|C90.31|ICD10CM|SOLITARY PLASMACYTOMA IN REMISSION|SOLITARY PLASMACYTOMA IN REMISSION
C4268569|T046|I97.821|ICD10CM|POSTPROCEDURAL CEREBROVASCULAR INFARCTION FOLLOWING OTHER SURGERY|POSTPROCEDURAL CEREBVASC INFARCTION FOLLOWING OTHER SURGERY
C4268568|T046|I97.820|ICD10CM|POSTPROCEDURAL CEREBROVASCULAR INFARCTION FOLLOWING CARDIAC SURGERY|POSTPROC CEREBVASC INFARCTION FOLLOWING CARDIAC SURGERY
C2891185|T037|T85.631A|ICD10CM|LEAKAGE OF INTRAPERITONEAL DIALYSIS CATHETER, INITIAL ENCOUNTER|LEAKAGE OF INTRAPERITONEAL DIALYSIS CATHETER, INIT ENCNTR
C2832594|T037|S06.821A|ICD10CM|INJURY OF LEFT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|INJ L INT CAROTID, INTCR W LOC OF 30 MINUTES OR LESS, INIT
C2891186|T037|T85.631D|ICD10CM|LEAKAGE OF INTRAPERITONEAL DIALYSIS CATHETER, SUBSEQUENT ENCOUNTER|LEAKAGE OF INTRAPERITONEAL DIALYSIS CATHETER, SUBS ENCNTR
C2889206|T047|M05.329|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP ELBOW
C2885173|T037|T61.782A|ICD10CM|OTHER SHELLFISH POISONING, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|OTH SHELLFISH POISONING, INTENTIONAL SELF-HARM, INIT ENCNTR
C2875142|T047|G40.911|ICD10CM|EPILEPSY, UNSPECIFIED, INTRACTABLE, WITH STATUS EPILEPTICUS|EPILEPSY, UNSPECIFIED, INTRACTABLE, WITH STATUS EPILEPTICUS
C2833174|T037|S12.031A|ICD10CM|NONDISPLACED POSTERIOR ARCH FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP POSTERIOR ARCH FX FIRST CERVCAL VERTEBRA, INIT
C2833175|T037|S12.031B|ICD10CM|NONDISPLACED POSTERIOR ARCH FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP POST ARCH FX FIRST CERVCAL VERTEBRA, INIT FOR OPN FX
C2875143|T047|G40.919|ICD10CM|EPILEPSY, UNSPECIFIED, INTRACTABLE, WITHOUT STATUS EPILEPTICUS|EPILEPSY, UNSP, INTRACTABLE, WITHOUT STATUS EPILEPTICUS
C2856967|T037|S72.062C|ICD10CM|DISPLACED ARTICULAR FRACTURE OF HEAD OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL ARTIC FX HEAD OF L FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2856966|T037|S72.062B|ICD10CM|DISPLACED ARTICULAR FRACTURE OF HEAD OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPLACED ARTIC FX HEAD OF L FEMUR, INIT FOR OPN FX TYPE I/2
C2856965|T037|S72.062A|ICD10CM|DISPLACED ARTICULAR FRACTURE OF HEAD OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED ARTICULAR FRACTURE OF HEAD OF LEFT FEMUR, INIT
C4237007|T048|F31.2|ICD10CM|BIPOLAR DISORDER, CURRENT EPISODE MANIC SEVERE WITH PSYCHOTIC FEATURES|BIPOLAR I DISORDER, CURRENT OR MOST RECENT EPISODE MANIC WITH PSYCHOTIC FEATURES
C2874872|T048|F31.0|ICD10CM|BIPOLAR DISORDER, CURRENT EPISODE HYPOMANIC|BIPOLAR DISORDER, CURRENT EPISODE HYPOMANIC
C2874885|T048|F31.4|ICD10CM|BIPOLAR DISORDER, CURRENT EPISODE DEPRESSED, SEVERE, WITHOUT PSYCHOTIC FEATURES|BIPOLAR DISORD, CRNT EPSD DEPRESS, SEV, W/O PSYCH FEATURES
C4237000|T048|F31.5|ICD10CM|BIPOLAR DISORDER, CURRENT EPISODE DEPRESSED, SEVERE, WITH PSYCHOTIC FEATURES|BIPOLAR I DISORDER, CURRENT OR MOST RECENT EPISODE DEPRESSED, WITH PSYCHOTIC FEATURES
C0005586|T048|F31|DMDICD10|BIPOLAR DISORDER, UNSPECIFIED|BIPOLARE AFFEKTIVE STOERUNG
C2901792|T047|M86.079|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED ANKLE AND FOOT|ACUTE HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED ANKLE AND FOOT
C2859971|T037|S78.011A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT RIGHT HIP JOINT, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION AT RIGHT HIP JOINT, INIT
C2901791|T047|M86.072|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, LEFT ANKLE AND FOOT|ACUTE HEMATOGENOUS OSTEOMYELITIS, LEFT ANKLE AND FOOT
C2901790|T047|M86.071|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, RIGHT ANKLE AND FOOT|ACUTE HEMATOGENOUS OSTEOMYELITIS, RIGHT ANKLE AND FOOT
C2873719|T191|D47.9|ICD10CM|NEOPLASM OF UNCERTAIN BEHAVIOR OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE, UNSPECIFIED|NEOPLM OF UNCRT BEHAV OF LYMPHOID,HEMATPOETC & REL TISS,UNSP
C2879542|T037|T46.6X2A|ICD10CM|POISONING BY ANTIHYPERLIPIDEMIC AND ANTIARTERIOSCLEROTIC DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY ANTIHYPERLIP AND ANTIARTERIO DRUGS, SELF-HARM, INIT
C2842084|T191|C50.111|ICD10CM|MALIGNANT NEOPLASM OF CENTRAL PORTION OF RIGHT FEMALE BREAST|MALIGNANT NEOPLASM OF CENTRAL PORTION OF RIGHT FEMALE BREAST
C2842085|T191|C50.112|ICD10CM|MALIGNANT NEOPLASM OF CENTRAL PORTION OF LEFT FEMALE BREAST|MALIGNANT NEOPLASM OF CENTRAL PORTION OF LEFT FEMALE BREAST
C1292778|T191|D47.1|DMDICD10|CHRONIC MYELOPROLIFERATIVE DISEASE|CHRONISCHE MYELOPROLIFERATIVE KRANKHEIT
C0040028|T047|D75.2|DMDICD10|ESSENTIAL (HEMORRHAGIC) THROMBOCYTHEMIA|ESSENTIELLE THROMBOZYTOSE
C0019068|T047|D76.2|DMDICD10|HEMOPHAGOCYTIC SYNDROME, INFECTION-ASSOCIATED|HAEMOPHAGOZYTAERES SYNDROM BEI INFEKTIONEN
C2873718|T191|D47.4|ICD10CM|OSTEOMYELOFIBROSIS|SECONDARY MYELOFIBROSIS IN MYELOPROLIFERATIVE DISEASE
C2890906|T037|T84.83XA|ICD10CM|HEMORRHAGE DUE TO INTERNAL ORTHOPEDIC PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|HEMORRHAGE DUE TO INTERNAL ORTHOPEDIC PROSTH DEV/GRFT, INIT
C2879544|T037|T46.6X2S|ICD10CM|POISONING BY ANTIHYPERLIPIDEMIC AND ANTIARTERIOSCLEROTIC DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY ANTIHYPERLIP AND ANTIARTERIO DRUGS, SLF-HRM, SQLA
C3264195|T047|H40.1214|ICD10CM|LOW-TENSION GLAUCOMA, RIGHT EYE, INDETERMINATE STAGE|LOW-TENSION GLAUCOMA, RIGHT EYE, INDETERMINATE STAGE
C3264192|T047|H40.1211|ICD10CM|LOW-TENSION GLAUCOMA, RIGHT EYE, MILD STAGE|LOW-TENSION GLAUCOMA, RIGHT EYE, MILD STAGE
C3264191|T047|H40.1210|ICD10CM|LOW-TENSION GLAUCOMA, RIGHT EYE, STAGE UNSPECIFIED|LOW-TENSION GLAUCOMA, RIGHT EYE, STAGE UNSPECIFIED
C3264194|T047|H40.1213|ICD10CM|LOW-TENSION GLAUCOMA, RIGHT EYE, SEVERE STAGE|LOW-TENSION GLAUCOMA, RIGHT EYE, SEVERE STAGE
C3264193|T047|H40.1212|ICD10CM|LOW-TENSION GLAUCOMA, RIGHT EYE, MODERATE STAGE|LOW-TENSION GLAUCOMA, RIGHT EYE, MODERATE STAGE
C0268558|T047|E72.50|ICD10CM|DISORDER OF GLYCINE METABOLISM, UNSPECIFIED|DISORDER OF GLYCINE METABOLISM, UNSPECIFIED
C0751748|T047||ICD10CM|NON-KETOTIC HYPERGLYCINEMIA
C0342739|T047|E72.52|ICD10CM|TRIMETHYLAMINURIA|TRIMETHYLAMINURIA
C1298681|T047|E72.53|ICD10CM|HYPEROXALURIA|OXALOSIS
C2874264|T047|E72.59|ICD10CM|OTHER DISORDERS OF GLYCINE METABOLISM|OTHER DISORDERS OF GLYCINE METABOLISM
C0343960|T047|B46.4|DMDICD10|DISSEMINATED MUCORMYCOSIS|DISSEMINIERTE MUKORMYKOSE
C0026718|T047|B46.5|DMDICD10|MUCORMYCOSIS, UNSPECIFIED|MUKORMYKOSE, NICHT NAEHER BEZEICHNET
C0339962|T047|B46.0|DMDICD10|PULMONARY MUCORMYCOSIS|MUKORMYKOSE DER LUNGE
C2882429|T047|I66.09|ICD10CM|OCCLUSION AND STENOSIS OF UNSPECIFIED MIDDLE CEREBRAL ARTERY|OCCLUSION AND STENOSIS OF UNSPECIFIED MIDDLE CEREBRAL ARTERY
C0348803|T047|B46.2|DMDICD10|GASTROINTESTINAL MUCORMYCOSIS|MUKORMYKOSE DES MAGEN-DARMTRAKTES
C2830240|T047|B46.3|ICD10CM|CUTANEOUS MUCORMYCOSIS|SUBCUTANEOUS MUCORMYCOSIS
C0839996|T047|M86.68|ICD10AM|OTHER CHRONIC OSTEOMYELITIS, OTHER SITE|OTHER CHRONIC OSTEOMYELITIS, OTHER SITE
C0839988|T047|M86.69|ICD10CM|OTHER CHRONIC OSTEOMYELITIS, MULTIPLE SITES|OTHER CHRONIC OSTEOMYELITIS, MULTIPLE SITES
C1396717|T047||ICD10CM|OTHER ZYGOMYCOSES
C2882426|T047|I66.01|ICD10CM|OCCLUSION AND STENOSIS OF RIGHT MIDDLE CEREBRAL ARTERY|OCCLUSION AND STENOSIS OF RIGHT MIDDLE CEREBRAL ARTERY
C2882427|T047|I66.02|ICD10CM|OCCLUSION AND STENOSIS OF LEFT MIDDLE CEREBRAL ARTERY|OCCLUSION AND STENOSIS OF LEFT MIDDLE CEREBRAL ARTERY
C2882428|T047|I66.03|ICD10CM|OCCLUSION AND STENOSIS OF BILATERAL MIDDLE CEREBRAL ARTERIES|OCCLUSION AND STENOSIS OF BILATERAL MIDDLE CEREBRAL ARTERIES
C2889214|T047|M05.341|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT HAND|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889215|T047|M05.342|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT HAND|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF LEFT HAND
C2889216|T047|M05.349|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP HAND
C4269552|T037|S02.671A|ICD10CM|FRACTURE OF ALVEOLUS OF RIGHT MANDIBLE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF ALVEOLUS OF RIGHT MANDIBLE, INIT
C2838683|T037|S34.125D|ICD10CM|INCOMPLETE LESION OF L5 LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|INCOMPLETE LESION OF L5 LEVEL OF LUMBAR SPINAL CORD, SUBS
C2838682|T037|S34.125A|ICD10CM|INCOMPLETE LESION OF L5 LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|INCOMPLETE LESION OF L5 LEVEL OF LUMBAR SPINAL CORD, INIT
C2878949|T037|T44.8X2S|ICD10CM|POISONING BY CENTRALLY-ACTING AND ADRENERGIC-NEURON-BLOCKING AGENTS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY CENTR-ACTING/ADREN-NEURN-BLOCK AGNT, SLF-HRM, SQLA
C2874563|T048|F13.950|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|SEDATV/HYP/ANXIOLYTC USE, UNSP W PSYCH DISORDER W DELUSIONS
C2874564|T048|F13.951|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|SEDATV/HYP/ANXIOLYTC USE, UNSP W PSYCH DISORDER W HALLUCIN
C2833958|T037|S14.131S|ICD10CM|ANTERIOR CORD SYNDROME AT C1 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|ANTERIOR CORD SYNDROME AT C1, SEQUELA
C4237407|T048|F13.959|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|SEDATIVE, HYPNOTIC, OR ANXIOLYTIC-INDUCED PSYCHOTIC DISORDER, WITHOUT USE DISORDER
C0020807|T047|J84.03|ICD10CM|IDIOPATHIC PULMONARY HEMOSIDEROSIS|ESSENTIAL BROWN INDURATION OF LUNG
C0155912|T047||ICD10CM|PULMONARY ALVEOLAR MICROLITHIASIS
C0034050|T047|J84.01|ICD10CM|ALVEOLAR PROTEINOSIS|ALVEOLAR PROTEINOSIS
C2833956|T037|S14.131A|ICD10CM|ANTERIOR CORD SYNDROME AT C1 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|ANTERIOR CORD SYNDROME AT C1, INIT
C3264392|T047|J84.09|ICD10CM|OTHER ALVEOLAR AND PARIETO-ALVEOLAR CONDITIONS|OTHER ALVEOLAR AND PARIETO-ALVEOLAR CONDITIONS
C2833957|T037|S14.131D|ICD10CM|ANTERIOR CORD SYNDROME AT C1 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|ANTERIOR CORD SYNDROME AT C1, SUBS
C2859140|T037|S73.001A|ICD10CM|UNSPECIFIED SUBLUXATION OF RIGHT HIP, INITIAL ENCOUNTER|UNSPECIFIED SUBLUXATION OF RIGHT HIP, INITIAL ENCOUNTER
C0265098|T190|I65.1|DMDICD10|OCCLUSION AND STENOSIS OF BASILAR ARTERY|VERSCHLUSS UND STENOSE DER A. BASILARIS
C4270126|T046|T82.818A|ICD10CM|EMBOLISM DUE TO VASCULAR PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|EMBOLISM DUE TO VASCULAR PROSTH DEV/GRFT, INITIAL ENCOUNTER
C0348637|T046|I65.8|DMDICD10|OCCLUSION AND STENOSIS OF OTHER PRECEREBRAL ARTERIES|VERSCHLUSS UND STENOSE SONSTIGER EXTRAKRANIELLER HIRNVERSORGENDER ARTERIE
C0155727|T047|I65.9|DMDICD10|OCCLUSION AND STENOSIS OF UNSPECIFIED PRECEREBRAL ARTERY|VERSCHLUSS UND STENOSE NICHT NAEHER BEZEICHNETER EXTRAKRANIELLER HIRNVERSORGENDER ARTERIE
C4270526|T046|T85.615A|ICD10CM|BREAKDOWN (MECHANICAL) OF OTHER NERVOUS SYSTEM DEVICE, IMPLANT OR GRAFT, INITIAL ENCOUNTER|BRKDWN OTHER NERVOUS SYS DEVICE, IMPLANT OR GRAFT, INIT
C2883255|T037|T48.992A|ICD10CM|POISONING BY OTHER AGENTS PRIMARILY ACTING ON THE RESPIRATORY SYSTEM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY OTH AGENTS PRIM ACT ON THE RESP SYS, SLF-HRM, INIT
C2855911|T037|S68.121S|ICD10CM|PARTIAL TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF LEFT INDEX FINGER, SEQUELA|PARTIAL TRAUMATIC MCP AMPUTATION OF L IDX FNGR, SEQUELA
C2890542|T037|T84.063A|ICD10CM|WEAR OF ARTICULAR BEARING SURFACE OF INTERNAL PROSTHETIC LEFT KNEE JOINT, INITIAL ENCOUNTER|WEAR OF ARTIC BEARING SURFACE OF INT PROSTH L KNEE JT, INIT
C2875372|T047|G90.519|ICD10CM|COMPLEX REGIONAL PAIN SYNDROME I OF UNSPECIFIED UPPER LIMB|COMPLEX REGIONAL PAIN SYNDROME I OF UNSPECIFIED UPPER LIMB
C2889962|T037|T82.391A|ICD10CM|OTHER MECHANICAL COMPLICATION OF CAROTID ARTERIAL GRAFT (BYPASS), INITIAL ENCOUNTER|MECH COMPL OF CAROTID ARTERIAL GRAFT (BYPASS), INIT ENCNTR
C2875369|T047|G90.511|ICD10CM|COMPLEX REGIONAL PAIN SYNDROME I OF RIGHT UPPER LIMB|COMPLEX REGIONAL PAIN SYNDROME I OF RIGHT UPPER LIMB
C2875370|T047|G90.512|ICD10CM|COMPLEX REGIONAL PAIN SYNDROME I OF LEFT UPPER LIMB|COMPLEX REGIONAL PAIN SYNDROME I OF LEFT UPPER LIMB
C2875371|T047|G90.513|ICD10CM|COMPLEX REGIONAL PAIN SYNDROME I OF UPPER LIMB, BILATERAL|COMPLEX REGIONAL PAIN SYNDROME I OF UPPER LIMB, BILATERAL
C2905756|T037|X78.1XXS|ICD10CM|INTENTIONAL SELF-HARM BY KNIFE, SEQUELA|INTENTIONAL SELF-HARM BY KNIFE, SEQUELA
C2900874|T046|M84.412A|ICD10CM|PATHOLOGICAL FRACTURE, LEFT SHOULDER, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, LEFT SHOULDER, INIT FOR FX
C2905755|T037|X78.1XXD|ICD10CM|INTENTIONAL SELF-HARM BY KNIFE, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY KNIFE, SUBSEQUENT ENCOUNTER
C2901935|T046|M87.00|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED BONE|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED BONE
C2905754|T037|X78.1XXA|ICD10CM|INTENTIONAL SELF-HARM BY KNIFE, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY KNIFE, INITIAL ENCOUNTER
C4509204|T046|I21.A9|ICD10CM|OTHER MYOCARDIAL INFARCTION TYPE|MYOCARDIAL INFARCTION ASSOCIATED WITH REVASCULARIZATION PROCEDURE
C2877922|T037|T41.202S|ICD10CM|POISONING BY UNSPECIFIED GENERAL ANESTHETICS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY UNSP GENERAL ANESTHETICS, SELF-HARM, SEQUELA
C2833841|T191|C06.80|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF UNSPECIFIED PARTS OF MOUTH|MALIGNANT NEOPLASM OF OVRLP SITES OF UNSP PARTS OF MOUTH
C2902423|T047|M90.50|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, UNSPECIFIED SITE|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, UNSP SITE
C2877252|T037|T38.892A|ICD10CM|POISONING BY OTHER HORMONES AND SYNTHETIC SUBSTITUTES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH HORMONES AND SYNTHETIC SUB, SELF-HARM, INIT
C2902452|T047||ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, OTHER SITE
C2902453|T047|M90.59|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, MULTIPLE SITES|OSTEONECROSIS IN DISEASES CLASSD ELSWHR, MULTIPLE SITES
C2877920|T037|T41.202A|ICD10CM|POISONING BY UNSPECIFIED GENERAL ANESTHETICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY UNSP GENERAL ANESTHETICS, SELF-HARM, INIT
C2890842|T037|T84.613A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL FIXATION DEVICE OF LEFT RADIUS, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INT FIX OF LEFT RADIUS, INIT
C2901082|T046|M84.474A|ICD10CM|PATHOLOGICAL FRACTURE, RIGHT FOOT, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, RIGHT FOOT, INIT ENCNTR FOR FRACTURE
C2900903|T046|M84.429A|ICD10CM|PATHOLOGICAL FRACTURE, UNSPECIFIED HUMERUS, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, UNSP HUMERUS, INIT FOR FX
C0275566|T047|A42.0|DMDICD10|PULMONARY ACTINOMYCOSIS|AKTINOMYKOSE DER LUNGE
C0349008|T047|A42.7|DMDICD10|ACTINOMYCOTIC SEPSIS|AKTINOMYKOTISCHE SEPSIS
C4521180|T047|I21.A1|ICD10CM|MYOCARDIAL INFARCTION TYPE 2|MYOCARDIAL INFARCTION TYPE 2
C2845942|T191|C74.02|ICD10CM|MALIGNANT NEOPLASM OF CORTEX OF LEFT ADRENAL GLAND|MALIGNANT NEOPLASM OF CORTEX OF LEFT ADRENAL GLAND
C2845941|T191|C74.01|ICD10CM|MALIGNANT NEOPLASM OF CORTEX OF RIGHT ADRENAL GLAND|MALIGNANT NEOPLASM OF CORTEX OF RIGHT ADRENAL GLAND
C2845940|T191|C74.00|ICD10CM|MALIGNANT NEOPLASM OF CORTEX OF UNSPECIFIED ADRENAL GLAND|MALIGNANT NEOPLASM OF CORTEX OF UNSPECIFIED ADRENAL GLAND
C2832049|T037|S06.2X9A|ICD10CM|DIFFUSE TRAUMATIC BRAIN INJURY WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|DIFFUSE TBI W LOSS OF CONSCIOUSNESS OF UNSP DURATION, INIT
C2835806|T037|S24.133D|ICD10CM|ANTERIOR CORD SYNDROME AT T7-T10 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|ANTERIOR CORD SYNDROME AT T7-T10, SUBS
C0478150|T184|R57.8|DMDICD10|OTHER SHOCK|SONSTIGE FORMEN DES SCHOCKS
C0036974|T046|R57.9|DMDICD10|SHOCK, UNSPECIFIED|SCHOCK, NICHT NAEHER BEZEICHNET
C2875333|T184||ICD10CM|SPASTIC HEMIPLEGIA AFFECTING LEFT NONDOMINANT SIDE
C2901588|T046|M84.68XA|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, OTHER SITE, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, OTH SITE, INIT FOR FX
C4270639|T046|T85.850A|ICD10CM|STENOSIS DUE TO NERVOUS SYSTEM PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|STENOSIS DUE TO NERVOUS SYSTEM PROSTH DEV/GRFT, INIT
C0154694|T047|G81.10|ICD10CM|SPASTIC HEMIPLEGIA AFFECTING UNSPECIFIED SIDE|SPASTIC HEMIPLEGIA AFFECTING UNSPECIFIED SIDE
C2875330|T184||ICD10CM|SPASTIC HEMIPLEGIA AFFECTING RIGHT DOMINANT SIDE
C2875331|T184||ICD10CM|SPASTIC HEMIPLEGIA AFFECTING LEFT DOMINANT SIDE
C2875332|T184||ICD10CM|SPASTIC HEMIPLEGIA AFFECTING RIGHT NONDOMINANT SIDE
C2889405|T047|M06.061|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, RIGHT KNEE|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, RIGHT KNEE
C2856082|T037|S68.629S|ICD10CM|PARTIAL TRAUMATIC TRANSPHALANGEAL AMPUTATION OF UNSPECIFIED FINGER, SEQUELA|PARTIAL TRAUMATIC TRNSPHAL AMP OF UNSP FINGER, SEQUELA
C2889406|T047|M06.062|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, LEFT KNEE|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, LEFT KNEE
C2835805|T037|S24.133A|ICD10CM|ANTERIOR CORD SYNDROME AT T7-T10 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|ANTERIOR CORD SYNDROME AT T7-T10, INIT
C4267900|T047|E08.3219|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|DIABETES WITH MILD NONP RTNOP WITH MACULAR EDEMA, UNSP
C2889407|T047|M06.06|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, UNSPECIFIED KNEE|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, KNEE
C4267898|T047|E08.3212|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|DIABETES WITH MILD NONP RTNOP WITH MACULAR EDEMA, LEFT EYE
C4267899|T047|E08.3213|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|DIABETES WITH MILD NONP RTNOP WITH MACULAR EDEMA, BILATERAL
C4267897|T047|E08.3211|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|DIABETES WITH MILD NONP RTNOP WITH MACULAR EDEMA, RIGHT EYE
C2874502|T048|F12.929|ICD10CM|CANNABIS USE, UNSPECIFIED WITH INTOXICATION, UNSPECIFIED|CANNABIS USE, UNSPECIFIED WITH INTOXICATION, UNSPECIFIED
C1401365|T047||ICD10CM|RICKETS, ACTIVE
C2874499|T048|F12.920|ICD10CM|CANNABIS USE, UNSPECIFIED WITH INTOXICATION, UNCOMPLICATED|CANNABIS USE, UNSPECIFIED WITH INTOXICATION, UNCOMPLICATED
C2874500|T048|F12.921|ICD10CM|CANNABIS USE, UNSPECIFIED WITH INTOXICATION DELIRIUM|CANNABIS USE, UNSPECIFIED WITH INTOXICATION DELIRIUM
C2874501|T048|F12.922|ICD10CM|CANNABIS USE, UNSPECIFIED WITH INTOXICATION WITH PERCEPTUAL DISTURBANCE|CANNABIS USE, UNSP W INTOXICATION W PERCEPTUAL DISTURBANCE
C2837590|T037|S32.040B|ICD10CM|WEDGE COMPRESSION FRACTURE OF FOURTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|WEDGE COMPRSN FX FOURTH LUM VERTEBRA, INIT FOR OPN FX
C2873947|T047|E08.9|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITHOUT COMPLICATIONS|DIABETES DUE TO UNDERLYING CONDITION W/O COMPLICATIONS
C2873946|T047|E08.8|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH UNSPECIFIED COMPLICATIONS|DIABETES DUE TO UNDERLYING CONDITION W UNSP COMPLICATIONS
C0153489|T191|C33|DMDICD10|MALIGNANT NEOPLASM OF TRACHEA|BOESARTIGE NEUBILDUNG DER TRACHEA
C2877764|T037|T40.7X2A|ICD10CM|POISONING BY CANNABIS (DERIVATIVES), INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY CANNABIS (DERIVATIVES), SELF-HARM, INIT
C1406705|T047||ICD10CM|TRIGEMINAL NEURALGIA
C0154729|T184|G50.1|DMDICD10|ATYPICAL FACIAL PAIN|ATYPISCHER GESICHTSSCHMERZ
C0477380|T047|G50.8|DMDICD10|OTHER DISORDERS OF TRIGEMINAL NERVE|SONSTIGE KRANKHEITEN DES N. TRIGEMINUS
C0152177|T047|G50|DMDICD10|DISORDER OF TRIGEMINAL NERVE, UNSPECIFIED|KRANKHEITEN DES N. TRIGEMINUS [V. HIRNNERV]
C2877766|T037|T40.7X2S|ICD10CM|POISONING BY CANNABIS (DERIVATIVES), INTENTIONAL SELF-HARM, SEQUELA|POISONING BY CANNABIS (DERIVATIVES), SELF-HARM, SEQUELA
C1955785|T047|I70.92|ICD10CM|CHRONIC TOTAL OCCLUSION OF ARTERY OF THE EXTREMITIES|TOTAL OCCLUSION OF ARTERY OF THE EXTREMITIES
C4269448|T037|S02.611B|ICD10CM|FRACTURE OF CONDYLAR PROCESS OF RIGHT MANDIBLE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF CONDYLAR PROCESS OF RIGHT MANDIBLE, 7THB
C4269447|T037|S02.611A|ICD10CM|FRACTURE OF CONDYLAR PROCESS OF RIGHT MANDIBLE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF CONDYLAR PROCESS OF RIGHT MANDIBLE, INIT
C0869206|T047|E88.2|DMDICD10|LIPOMATOSIS, NOT ELSEWHERE CLASSIFIED|LIPOMATOSE, ANDERENORTS NICHT KLASSIFIZIERT
C2856099|T037|S68.721A|ICD10CM|PARTIAL TRAUMATIC TRANSMETACARPAL AMPUTATION OF RIGHT HAND, INITIAL ENCOUNTER|PARTIAL TRAUMATIC TRANSMETCRPL AMP OF RIGHT HAND, INIT
C2861681|T191|D03.71|ICD10CM|MELANOMA IN SITU OF RIGHT LOWER LIMB, INCLUDING HIP|MELANOMA IN SITU OF RIGHT LOWER LIMB, INCLUDING HIP
C2861680|T191|D03.70|ICD10CM|MELANOMA IN SITU OF UNSPECIFIED LOWER LIMB, INCLUDING HIP|MELANOMA IN SITU OF UNSPECIFIED LOWER LIMB, INCLUDING HIP
C2856101|T037|S68.721S|ICD10CM|PARTIAL TRAUMATIC TRANSMETACARPAL AMPUTATION OF RIGHT HAND, SEQUELA|PARTIAL TRAUMATIC TRANSMETCRPL AMP OF RIGHT HAND, SEQUELA
C2831986|T037|S06.1X3S|ICD10CM|TRAUMATIC CEREBRAL EDEMA WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, SEQUELA|TRAUMATIC CEREBRAL EDEMA W LOC OF 1-5 HRS 59 MIN, SEQUELA
C2882374|T047|I63.339|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF UNSPECIFIED POSTERIOR CEREBRAL ARTERY|CEREBRAL INFRC DUE TO THOMBOS UNSP POSTERIOR CEREBRAL ARTERY
C2831938|T037|S06.0X1S|ICD10CM|CONCUSSION WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|CONCUSSION W LOC OF 30 MINUTES OR LESS, SEQUELA
C2873912|T047|E08.36|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH DIABETIC CATARACT|DIABETES DUE TO UNDERLYING CONDITION W DIABETIC CATARACT
C2873913|T047|E08.39|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH OTHER DIABETIC OPHTHALMIC COMPLICATION|DIABETES DUE TO UNDRL CONDITION W OTH DIABETIC OPTH COMP
C2905738|T037|X77.3XXA|ICD10CM|INTENTIONAL SELF-HARM BY HOT HOUSEHOLD APPLIANCES, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY HOT HOUSEHOLD APPLIANCES, INIT
C2905739|T037|X77.3XXD|ICD10CM|INTENTIONAL SELF-HARM BY HOT HOUSEHOLD APPLIANCES, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY HOT HOUSEHOLD APPLIANCES, SUBS
C2882372|T047|I63.331|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF RIGHT POSTERIOR CEREBRAL ARTERY|CEREBRAL INFRC DUE TO THOMBOS OF RIGHT POST CEREBRAL ARTERY
C0342181|T046||ICD10CM|OTHER SPECIFIED DISORDERS OF THYROID
C4268483|T047|I63.333|ICD10CM|CEREBRAL INFARCTION TO THROMBOSIS OF BILATERAL POSTERIOR CEREBRAL ARTERIES|CEREBRAL INFRC TO THOMBOS OF BI POSTERIOR CEREBRAL ARTERIES
C2831984|T037|S06.1X3A|ICD10CM|TRAUMATIC CEREBRAL EDEMA WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|TRAUMATIC CEREBRAL EDEMA W LOC OF 1-5 HRS 59 MIN, INIT
C2842104|T191|C50.329|ICD10CM|MALIGNANT NEOPLASM OF LOWER-INNER QUADRANT OF UNSPECIFIED MALE BREAST|MALIG NEOPLASM OF LOWER-INNER QUADRANT OF UNSP MALE BREAST
C2842103|T191|C50.322|ICD10CM|MALIGNANT NEOPLASM OF LOWER-INNER QUADRANT OF LEFT MALE BREAST|MALIG NEOPLASM OF LOWER-INNER QUADRANT OF LEFT MALE BREAST
C2842102|T191|C50.321|ICD10CM|MALIGNANT NEOPLASM OF LOWER-INNER QUADRANT OF RIGHT MALE BREAST|MALIG NEOPLASM OF LOWER-INNER QUADRANT OF RIGHT MALE BREAST
C2905740|T037|X77.3XXS|ICD10CM|INTENTIONAL SELF-HARM BY HOT HOUSEHOLD APPLIANCES, SEQUELA|INTENTIONAL SELF-HARM BY HOT HOUSEHOLD APPLIANCES, SEQUELA
C2884945|T037|T59.7X2A|ICD10CM|TOXIC EFFECT OF CARBON DIOXIDE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CARBON DIOXIDE, INTENTIONAL SELF-HARM, INIT
C4268145|T047|E13.3491|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|OTH DIAB WITH SEVERE NONP RTNOP WITHOUT MACULAR EDEMA, R EYE
C4268146|T047|E13.3492|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|OTH DIAB WITH SEVERE NONP RTNOP WITHOUT MACULAR EDEMA, L EYE
C4268147|T047|E13.3493|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|OTH DIAB WITH SEVERE NONP RTNOP WITHOUT MACULAR EDEMA, BI
C0242006|T047||ICD10CM|MYELOFIBROSIS
C4268148|T047|E13.3499|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|OTH DIAB WITH SEVERE NONP RTNOP WITHOUT MACULAR EDEMA, UNSP
C2857207|T037|S72.114C|ICD10CM|NONDISPLACED FRACTURE OF GREATER TROCHANTER OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF GREATER TROCHANTER OF R FEMR, 7THC
C0272285|T047|D75.82|ICD10CM|HEPARIN INDUCED THROMBOCYTOPENIA (HIT)|HEPARIN INDUCED THROMBOCYTOPENIA (HIT)
C2833896|T037|S14.114S|ICD10CM|COMPLETE LESION AT C4 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|COMPLETE LESION AT C4 LEVEL OF CERVICAL SPINAL CORD, SEQUELA
C2887220|T047|I83.219|ICD10CM|VARICOSE VEINS OF RIGHT LOWER EXTREMITY WITH BOTH ULCER OF UNSPECIFIED SITE AND INFLAMMATION|VARICOS VN OF R LOW EXTREM W ULC OF UNSP SITE AND INFLAM
C2887219|T047|I83.218|ICD10CM|VARICOSE VEINS OF RIGHT LOWER EXTREMITY WITH BOTH ULCER OF OTHER PART OF LOWER EXTREMITY AND INFLAMMATION|VARICOS VN OF R LOW EXTREM W ULC OTH PRT LOW EXTRM & INFLAM
C2887212|T047|I83.211|ICD10CM|VARICOSE VEINS OF RIGHT LOWER EXTREMITY WITH BOTH ULCER OF THIGH AND INFLAMMATION|VARICOS VN OF R LOW EXTREM W ULC OF THIGH AND INFLAMMATION
C2833895|T037|S14.114D|ICD10CM|COMPLETE LESION AT C4 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|COMPLETE LESION AT C4 LEVEL OF CERVICAL SPINAL CORD, SUBS
C2887214|T047|I83.213|ICD10CM|VARICOSE VEINS OF RIGHT LOWER EXTREMITY WITH BOTH ULCER OF ANKLE AND INFLAMMATION|VARICOS VN OF R LOW EXTREM W ULC OF ANKLE AND INFLAMMATION
C2887213|T047|I83.212|ICD10CM|VARICOSE VEINS OF RIGHT LOWER EXTREMITY WITH BOTH ULCER OF CALF AND INFLAMMATION|VARICOS VN OF R LOW EXTREM W ULC OF CALF AND INFLAMMATION
C2887218|T047|I83.215|ICD10CM|VARICOSE VEINS OF RIGHT LOWER EXTREMITY WITH BOTH ULCER OTHER PART OF FOOT AND INFLAMMATION|VARICOS VN OF R LOW EXTREM W ULC OTH PART OF FOOT AND INFLAM
C2887216|T047|I83.214|ICD10CM|VARICOSE VEINS OF RIGHT LOWER EXTREMITY WITH BOTH ULCER OF HEEL AND MIDFOOT AND INFLAMMATION|VARICOS VN OF R LOW EXTREM W ULC OF HEEL & MIDFT AND INFLAM
C0010823|T047|B25.9|DMDICD10|CYTOMEGALOVIRAL DISEASE, UNSPECIFIED|ZYTOMEGALIE, NICHT NAEHER BEZEICHNET
C0348218|T047|B25.8|DMDICD10|OTHER CYTOMEGALOVIRAL DISEASES|SONSTIGE ZYTOMEGALIE
C2869847|T037|S98.221A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF TWO OR MORE RIGHT LESSER TOES, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP OF TWO OR MORE RIGHT LESSER TOES, INIT
C2869848|T037|S98.221D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF TWO OR MORE RIGHT LESSER TOES, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMP OF TWO OR MORE RIGHT LESSER TOES, SUBS
C0341465|T047|B25.2|DMDICD10|CYTOMEGALOVIRAL PANCREATITIS|PANKREATITIS DURCH ZYTOMEGALIEVIREN
C0276252|T047|B25.1|DMDICD10|CYTOMEGALOVIRAL HEPATITIS|HEPATITIS DURCH ZYTOMEGALIEVIREN
C0276253|T047|B25.0|DMDICD10|CYTOMEGALOVIRAL PNEUMONITIS|PNEUMONIE DURCH ZYTOMEGALIEVIREN
C2901364|T046|M84.60XA|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, UNSPECIFIED SITE, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, UNSP SITE, INIT FOR FX
C2874382|T048|F10.19|ICD10CM|ALCOHOL ABUSE WITH UNSPECIFIED ALCOHOL-INDUCED DISORDER|ALCOHOL ABUSE WITH UNSPECIFIED ALCOHOL-INDUCED DISORDER
C2869849|T037|S98.221S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF TWO OR MORE RIGHT LESSER TOES, SEQUELA|PARTIAL TRAUM AMP OF TWO OR MORE RIGHT LESSER TOES, SEQUELA
C4268203|T048|F10.14|ICD10CM|ALCOHOL ABUSE WITH ALCOHOL-INDUCED MOOD DISORDER|ALCOHOL USE DISORDER, MILD, WITH ALCOHOL-INDUCED DEPRESSIVE DISORDER
C2905780|T037|X81.0XXS|ICD10CM|INTENTIONAL SELF-HARM BY JUMPING OR LYING IN FRONT OF MOTOR VEHICLE, SEQUELA|SELF-HARM BY JUMPING OR LYING IN FRONT OF MTR VEH, SEQUELA
C2832282|T037|S06.355A|ICD10CM|TRAUMATIC HEMORRHAGE OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, INITIAL ENCOUNTER|TRAUM HEMOR LEFT CEREBRUM W LOC >24 HR W RET CONSC LEV, INIT
C2901829|T047|M86.241|ICD10CM|SUBACUTE OSTEOMYELITIS, RIGHT HAND|SUBACUTE OSTEOMYELITIS, RIGHT HAND
C2905779|T037|X81.0XXD|ICD10CM|INTENTIONAL SELF-HARM BY JUMPING OR LYING IN FRONT OF MOTOR VEHICLE, SUBSEQUENT ENCOUNTER|SELF-HARM BY JUMPING OR LYING IN FRONT OF MTR VEH, SUBS
C2901830|T047|M86.242|ICD10CM|SUBACUTE OSTEOMYELITIS, LEFT HAND|SUBACUTE OSTEOMYELITIS, LEFT HAND
C2911419|T033|Z89.442|ICD10CM|ACQUIRED ABSENCE OF LEFT ANKLE|ACQUIRED ABSENCE OF LEFT ANKLE
C1260398|T047|D57.219|ICD10CM|SICKLE-CELL/HB-C DISEASE WITH CRISIS, UNSPECIFIED|SICKLE-CELL/HB-C DISEASE WITH CRISIS, UNSPECIFIED
C2905778|T037|X81.0XXA|ICD10CM|INTENTIONAL SELF-HARM BY JUMPING OR LYING IN FRONT OF MOTOR VEHICLE, INITIAL ENCOUNTER|SELF-HARM BY JUMPING OR LYING IN FRONT OF MTR VEH, INIT
C0236764|T048|F33.41|ICD10CM|MAJOR DEPRESSIVE DISORDER, RECURRENT, IN PARTIAL REMISSION|MAJOR DEPRESSIVE DISORDER, RECURRENT, IN PARTIAL REMISSION
C2874933|T048|F33.4|ICD10CM|MAJOR DEPRESSIVE DISORDER, RECURRENT, IN REMISSION, UNSPECIFIED|MAJOR DEPRESSIVE DISORDER, RECURRENT, IN REMISSION
C2891329|T037|T87.40|ICD10CM|INFECTION OF AMPUTATION STUMP, UNSPECIFIED EXTREMITY|INFECTION OF AMPUTATION STUMP, UNSPECIFIED EXTREMITY
C3665667|T048|F33.42|ICD10CM|MAJOR DEPRESSIVE DISORDER, RECURRENT, IN FULL REMISSION|MAJOR DEPRESSIVE DISORDER, RECURRENT, IN FULL REMISSION
C2873764|T047||ICD10CM|SICKLE-CELL/HB-C DISEASE WITH SPLENIC SEQUESTRATION
C2873763|T047||ICD10CM|SICKLE-CELL/HB-C DISEASE WITH ACUTE CHEST SYNDROME
C2882263|T046|I46.2|ICD10CM|CARDIAC ARREST DUE TO UNDERLYING CARDIAC CONDITION|CARDIAC ARREST DUE TO UNDERLYING CARDIAC CONDITION
C2905762|T037|X78.8XXA|ICD10CM|INTENTIONAL SELF-HARM BY OTHER SHARP OBJECT, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY OTHER SHARP OBJECT, INIT ENCNTR
C2882265|T046|I46.9|ICD10CM|CARDIAC ARREST, CAUSE UNSPECIFIED|CARDIAC ARREST, CAUSE UNSPECIFIED
C2882264|T046|I46.8|ICD10CM|CARDIAC ARREST DUE TO OTHER UNDERLYING CONDITION|CARDIAC ARREST DUE TO OTHER UNDERLYING CONDITION
C2905763|T037|X78.8XXD|ICD10CM|INTENTIONAL SELF-HARM BY OTHER SHARP OBJECT, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY OTHER SHARP OBJECT, SUBS ENCNTR
C4270284|T046|T83.25XA|ICD10CM|EXPOSURE OF GRAFT OF URINARY ORGAN, INITIAL ENCOUNTER|EXPOSURE OF GRAFT OF URINARY ORGAN, INITIAL ENCOUNTER
C2905764|T037|X78.8XXS|ICD10CM|INTENTIONAL SELF-HARM BY OTHER SHARP OBJECT, SEQUELA|INTENTIONAL SELF-HARM BY OTHER SHARP OBJECT, SEQUELA
C2881302|T047|H49.812|ICD10CM|KEARNS-SAYRE SYNDROME, LEFT EYE|KEARNS-SAYRE SYNDROME, LEFT EYE
C2881303|T047|H49.813|ICD10CM|KEARNS-SAYRE SYNDROME, BILATERAL|KEARNS-SAYRE SYNDROME, BILATERAL
C2881301|T047|H49.811|ICD10CM|KEARNS-SAYRE SYNDROME, RIGHT EYE|KEARNS-SAYRE SYNDROME, RIGHT EYE
C2842031|T191|C47.12|ICD10CM|MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF LEFT UPPER LIMB, INCLUDING SHOULDER|MALIG NEOPLM OF PRPH NERVES OF LEFT UPPER LIMB, INC SHOULDER
C2842029|T191|C47.10|ICD10CM|MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF UNSPECIFIED UPPER LIMB, INCLUDING SHOULDER|MALIG NEOPLM OF PRPH NERVES OF UNSP UPPER LIMB, INC SHOULDER
C2842030|T191|C47.11|ICD10CM|MALIGNANT NEOPLASM OF PERIPHERAL NERVES OF RIGHT UPPER LIMB, INCLUDING SHOULDER|MALIG NEOPLM OF PRPH NERVES OF RIGHT UPPER LIMB, INC SHLDR
C2874747|T048||ICD10CM|INHALANT ABUSE WITH INTOXICATION, UNCOMPLICATED
C2881304|T047|H49.819|ICD10CM|KEARNS-SAYRE SYNDROME, UNSPECIFIED EYE|KEARNS-SAYRE SYNDROME, UNSPECIFIED EYE
C2890011|T037|T82.513A|ICD10CM|BREAKDOWN (MECHANICAL) OF BALLOON (COUNTERPULSATION) DEVICE, INITIAL ENCOUNTER|BREAKDOWN OF BALLOON (COUNTERPULSATION) DEVICE, INIT
C2889598|T047|M08.48|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, VERTEBRAE|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, VERTEBRAE
C0837721|T047|M08.40|ICD10AM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED SITE|PAUCIARTICULAR JUVENILE ARTHRITIS, MULTIPLE SITES
C2888661|T047|L97.204|ICD10CM|NON-PRESSURE CHRONIC ULCER OF UNSPECIFIED CALF WITH NECROSIS OF BONE|NON-PRESSURE CHRONIC ULCER OF UNSP CALF W NECROSIS OF BONE
C0348653|T047|I79.1|DMDICD10|AORTITIS IN DISEASES CLASSIFIED ELSEWHERE|AORTITIS BEI ANDERENORTS KLASSIFIZIERTEN KRANKHEITEN
C0348652|T190|I79.0|DMDICD10|ANEURYSM OF AORTA IN DISEASES CLASSIFIED ELSEWHERE|AORTENANEURYSMA BEI ANDERENORTS KLASSIFIZIERTEN KRANKHEITEN
C2889579|T047|M08.422|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, LEFT ELBOW|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, LEFT ELBOW
C2889578|T047|M08.421|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, RIGHT ELBOW|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, RIGHT ELBOW
C0348654|T047|I79.8|DMDICD10|OTHER DISORDERS OF ARTERIES, ARTERIOLES AND CAPILLARIES IN DISEASES CLASSIFIED ELSEWHERE|SONSTIGE KRANKHEITEN DER ARTERIEN, ARTERIOLEN UND KAPILLAREN BEI ANDERENORTS KLASSIFIZIERTEN KRANKHEITEN
C2889580|T047|M08.429|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED ELBOW|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED ELBOW
C0264444|T047|J63.5|DMDICD10|STANNOSIS|STANNOSE
C0037061|T047|J63.4|DMDICD10|SIDEROSIS|SIDEROSE
C0348695|T047|J63.6|ICD10CM|PNEUMOCONIOSIS DUE TO OTHER SPECIFIED INORGANIC DUSTS|PNEUMOCONIOSIS DUE TO OTHER SPECIFIED INORGANIC DUSTS
C0264437|T047|J63.1|DMDICD10|BAUXITE FIBROSIS (OF LUNG)|BAUXITFIBROSE (LUNGE)
C0311227|T047|J63.0|DMDICD10|ALUMINOSIS (OF LUNG)|ALUMINOSE (LUNGE)
C0264439|T047|J63.3|DMDICD10|GRAPHITE FIBROSIS (OF LUNG)|GRAPHITFIBROSE (LUNGE)
C0494309|T046|E23.1|DMDICD10|DRUG-INDUCED HYPOPITUITARISM|ARZNEIMITTELINDUZIERTER HYPOPITUITARISMUS
C2837632|T037|S32.051A|ICD10CM|STABLE BURST FRACTURE OF FIFTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|STABLE BURST FRACTURE OF FIFTH LUMBAR VERTEBRA, INIT
C2837633|T037|S32.051B|ICD10CM|STABLE BURST FRACTURE OF FIFTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|STABLE BURST FRACTURE OF FIFTH LUM VERTEBRA, INIT FOR OPN FX
C2902441|T047|M90.551|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, RIGHT THIGH|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, RIGHT THIGH
C2877893|T037|T41.1X2A|ICD10CM|POISONING BY INTRAVENOUS ANESTHETICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY INTRAVENOUS ANESTHETICS, SELF-HARM, INIT
C2890055|T037|T82.528A|ICD10CM|DISPLACEMENT OF OTHER CARDIAC AND VASCULAR DEVICES AND IMPLANTS, INITIAL ENCOUNTER|DISPLACMNT OF CARDIAC AND VASCULAR DEVICES AND IMPLNT, INIT
C2832301|T037|S06.359S|ICD10CM|TRAUMATIC HEMORRHAGE OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|TRAUM HEMOR LEFT CEREBRUM W LOC OF UNSP DURATION, SEQUELA
C2873842|T047|D80.0|ICD10CM|HEREDITARY HYPOGAMMAGLOBULINEMIA|X-LINKED AGAMMAGLOBULINEMIA [BRUTON] (WITH GROWTH HORMONE DEFICIENCY)
C2873843|T047|D80.1|ICD10CM|NONFAMILIAL HYPOGAMMAGLOBULINEMIA|COMMON VARIABLE AGAMMAGLOBULINEMIA [CVAGAMMA]
C4049006|T047|D80.2|DMDICD10|SELECTIVE DEFICIENCY OF IMMUNOGLOBULIN A [IGA]|SELEKTIVER IMMUNGLOBULIN-A-MANGEL [IGA-MANGEL]
C0162539|T047|D80.3|DMDICD10|SELECTIVE DEFICIENCY OF IMMUNOGLOBULIN G [IGG] SUBCLASSES|SELEKTIVER MANGEL AN IMMUNGLOBULIN-G-SUBKLASSEN [IGG-SUBKLASSEN]
C2887842|T047|K51.913|ICD10CM|ULCERATIVE COLITIS, UNSPECIFIED WITH FISTULA|ULCERATIVE COLITIS, UNSPECIFIED WITH FISTULA
C0740331|T047|D80.5|DMDICD10|IMMUNODEFICIENCY WITH INCREASED IMMUNOGLOBULIN M [IGM]|IMMUNDEFEKT BEI ERHOEHTEM IMMUNGLOBULIN M [IGM]
C2887840|T047|K51.911|ICD10CM|ULCERATIVE COLITIS, UNSPECIFIED WITH RECTAL BLEEDING|ULCERATIVE COLITIS, UNSPECIFIED WITH RECTAL BLEEDING
C0272238|T047|D80.7|DMDICD10|TRANSIENT HYPOGAMMAGLOBULINEMIA OF INFANCY|TRANSITORISCHE HYPOGAMMAGLOBULINAEMIE IM KINDESALTER
C3248381|T047|D80.8|ICD10CM|OTHER IMMUNODEFICIENCIES WITH PREDOMINANTLY ANTIBODY DEFECTS|KAPPA LIGHT CHAIN DEFICIENCY
C0494248|T047|D80|DMDICD10|IMMUNODEFICIENCY WITH PREDOMINANTLY ANTIBODY DEFECTS, UNSPECIFIED|IMMUNDEFEKT MIT VORHERRSCHENDEM ANTIKOERPERMANGEL
C4269398|T037|S02.40DA|ICD10CM|MAXILLARY FRACTURE, LEFT SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|MAXILLARY FRACTURE, LEFT SIDE, INIT
C0153645|T191|C70.0|DMDICD10|MALIGNANT NEOPLASM OF CEREBRAL MENINGES|BOESARTIGE NEUBILDUNG: HIRNHAEUTE
C2887845|T047|K51.919|ICD10CM|ULCERATIVE COLITIS, UNSPECIFIED WITH UNSPECIFIED COMPLICATIONS|ULCERATIVE COLITIS, UNSP WITH UNSPECIFIED COMPLICATIONS
C2887844|T047|K51.918|ICD10CM|ULCERATIVE COLITIS, UNSPECIFIED WITH OTHER COMPLICATION|ULCERATIVE COLITIS, UNSPECIFIED WITH OTHER COMPLICATION
C2883684|T037|T50.6X2A|ICD10CM|POISONING BY ANTIDOTES AND CHELATING AGENTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ANTIDOTES AND CHELATING AGENTS, SELF-HARM, INIT
C2890600|T037|T84.115A|ICD10CM|BREAKDOWN (MECHANICAL) OF INTERNAL FIXATION DEVICE OF LEFT FEMUR, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF INT FIX OF LEFT FEMUR, INIT
C2883686|T037|T50.6X2S|ICD10CM|POISONING BY ANTIDOTES AND CHELATING AGENTS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY ANTIDOTES AND CHELATING AGENTS, SELF-HARM, SEQUELA
C2832184|T037|S06.331S|ICD10CM|CONTUSION AND LACERATION OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|CONTUS/LAC CEREB, W LOC OF 30 MINUTES OR LESS, SEQUELA
C2890222|T037|T83.030A|ICD10CM|LEAKAGE OF CYSTOSTOMY CATHETER, INITIAL ENCOUNTER|LEAKAGE OF CYSTOSTOMY CATHETER, INITIAL ENCOUNTER
C2835198|T037|S22.011B|ICD10CM|STABLE BURST FRACTURE OF FIRST THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|STABLE BURST FX FIRST THOR VERTEBRA, INIT FOR OPN FX
C2835197|T037|S22.011A|ICD10CM|STABLE BURST FRACTURE OF FIRST THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|STABLE BURST FRACTURE OF FIRST THORACIC VERTEBRA, INIT
C2832182|T037|S06.331A|ICD10CM|CONTUSION AND LACERATION OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|CONTUS/LAC CEREB, W LOC OF 30 MINUTES OR LESS, INIT
C3263995|T047|G40.A19|ICD10CM|ABSENCE EPILEPTIC SYNDROME, INTRACTABLE, WITHOUT STATUS EPILEPTICUS|ABSENCE EPILEPTIC SYNDROME, INTRACTABLE, W/O STAT EPI
C2837604|T037|S32.042B|ICD10CM|UNSTABLE BURST FRACTURE OF FOURTH LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSTABLE BURST FX FOURTH LUM VERTEBRA, INIT FOR OPN FX
C3263994|T047|G40.A11|ICD10CM|ABSENCE EPILEPTIC SYNDROME, INTRACTABLE, WITH STATUS EPILEPTICUS|ABSENCE EPILEPTIC SYNDROME, INTRACTABLE, W STAT EPI
C4268013|T047|E10.3213|ICD10CM|TYPE 1 DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|TYPE 1 DIABETES WITH MILD NONP RTNOP WITH MACULAR EDEMA, BI
C4268012|T047|E10.3212|ICD10CM|TYPE 1 DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|TYPE 1 DIAB WITH MILD NONP RTNOP WITH MACULAR EDEMA, L EYE
C4270423|T046|T83.79XA|ICD10CM|OTHER SPECIFIED COMPLICATIONS DUE TO OTHER GENITOURINARY PROSTHETIC MATERIALS, INITIAL ENCOUNTER|OTH COMP DUE TO OTHER GU PROSTHETIC MATERIALS, INIT
C4267969|T047|E09.3399|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|DRUG/CHEM DIAB WITH MOD NONP RTNOP WITHOUT MCLR EDEMA, UNSP
C4267967|T047|E09.3392|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|DRUG/CHEM DIAB WITH MOD NONP RTNOP WITHOUT MCLR EDEMA, L EYE
C4267968|T047|E09.3393|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|DRUG/CHEM DIAB WITH MOD NONP RTNOP WITHOUT MACULAR EDEMA, BI
C4267966|T047|E09.3391|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH MODERATE NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|DRUG/CHEM DIAB WITH MOD NONP RTNOP WITHOUT MCLR EDEMA, R EYE
C0347054|T191|C77.3|ICD10CM|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF AXILLA AND UPPER LIMB LYMPH NODES|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF PECTORAL LYMPH NODES
C0686655|T191|C77.2|DMDICD10|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF INTRA-ABDOMINAL LYMPH NODES|SEKUNDAERE UND NICHT NAEHER BEZEICHNETE BOESARTIGE NEUBILDUNG: INTRAABDOMINALE LYMPHKNOTEN
C0686645|T191|C77.1|DMDICD10|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF INTRATHORACIC LYMPH NODES|SEKUNDAERE UND NICHT NAEHER BEZEICHNETE BOESARTIGE NEUBILDUNG: INTRATHORAKALE LYMPHKNOTEN
C0864998|T191|C77.0|ICD10CM|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF LYMPH NODES OF HEAD, FACE AND NECK|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF SUPRACLAVICULAR LYMPH NODES
C0686689|T191|C77.5|DMDICD10|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF INTRAPELVIC LYMPH NODES|SEKUNDAERE UND NICHT NAEHER BEZEICHNETE BOESARTIGE NEUBILDUNG: INTRAPELVINE LYMPHKNOTEN
C0347055|T191|C77.4|DMDICD10|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF INGUINAL AND LOWER LIMB LYMPH NODES|SEKUNDAERE UND NICHT NAEHER BEZEICHNETE BOESARTIGE NEUBILDUNG: INGUINALE LYMPHKNOTEN UND LYMPHKNOTEN DER UNTEREN EXTREMITAET
C0686619|T191|C77.9|DMDICD10|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF LYMPH NODE, UNSPECIFIED|SEKUNDAERE UND NICHT NAEHER BEZEICHNETE BOESARTIGE NEUBILDUNG: LYMPHKNOTEN, NICHT NAEHER BEZEICHNET
C0348382|T191|C77.8|DMDICD10|SECONDARY AND UNSPECIFIED MALIGNANT NEOPLASM OF LYMPH NODES OF MULTIPLE REGIONS|SEKUNDAERE UND NICHT NAEHER BEZEICHNETE BOESARTIGE NEUBILDUNG: LYMPHKNOTEN MEHRERER REGIONEN
C2884170|T037|T52.8X2S|ICD10CM|TOXIC EFFECT OF OTHER ORGANIC SOLVENTS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF ORGANIC SOLVENTS, SELF-HARM, SEQUELA
C2890723|T037|T84.228A|ICD10CM|DISPLACEMENT OF INTERNAL FIXATION DEVICE OF OTHER BONES, INITIAL ENCOUNTER|DISPLACEMENT OF INTERNAL FIXATION DEVICE OF OTH BONES, INIT
C2856861|T037|S72.045A|ICD10CM|NONDISPLACED FRACTURE OF BASE OF NECK OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF BASE OF NECK OF LEFT FEMUR, INIT FOR CLOS FX
C0400883|T047|K55|DMDICD10|VASCULAR DISORDER OF INTESTINE, UNSPECIFIED|GEFAESSKRANKHEITEN DES DARMES
C0348740|T047|K55.8|DMDICD10|OTHER VASCULAR DISORDERS OF INTESTINE|SONSTIGE GEFAESSKRANKHEITEN DES DARMES
C2859063|T037|S72.8X9C|ICD10CM|OTHER FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|OTH FRACTURE OF UNSP FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C1412000|T047|K55.1|ICD10CM|CHRONIC VASCULAR DISORDERS OF INTESTINE|MESENTERIC VASCULAR INSUFFICIENCY
C2857942|T037|S72.342A|ICD10CM|DISPLACED SPIRAL FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED SPIRAL FRACTURE OF SHAFT OF LEFT FEMUR, INIT
C2857943|T037|S72.342B|ICD10CM|DISPLACED SPIRAL FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL SPIRAL FX SHAFT OF L FEMUR, INIT FOR OPN FX TYPE I/2
C2857944|T037|S72.342C|ICD10CM|DISPLACED SPIRAL FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL SPIRAL FX SHAFT OF L FEMR, INIT FOR OPN FX TYPE 3A/B/C
C2889302|T047|M05.622|ICD10CM|RHEUMATOID ARTHRITIS OF LEFT ELBOW WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF L ELBOW W INVOLV OF ORGANS AND SYSTEMS
C2889153|T047|M05.151|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT HIP|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889154|T047|M05.152|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT HIP|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT HIP
C2889301|T047|M05.621|ICD10CM|RHEUMATOID ARTHRITIS OF RIGHT ELBOW WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF R ELBOW W INVOLV OF ORGANS AND SYSTEMS
C2889152|T047|M05.159|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP
C2856930|T037|S72.059A|ICD10CM|UNSPECIFIED FRACTURE OF HEAD OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF HEAD OF UNSP FEMUR, INIT FOR CLOS FX
C2889303|T047|M05.629|ICD10CM|RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF UNSP ELBOW W INVOLV OF ORGANS AND SYSTEMS
C2842055|T191|C4A.21|ICD10CM|MERKEL CELL CARCINOMA OF RIGHT EAR AND EXTERNAL AURICULAR CANAL|MERKEL CELL CARCINOMA OF RIGHT EAR AND EXTERNAL AURIC CANAL
C2977924|T191|C4A.20|ICD10CM|MERKEL CELL CARCINOMA OF UNSPECIFIED EAR AND EXTERNAL AURICULAR CANAL|MERKEL CELL CARCINOMA OF UNSP EAR AND EXTERNAL AURIC CANAL
C2842056|T191|C4A.22|ICD10CM|MERKEL CELL CARCINOMA OF LEFT EAR AND EXTERNAL AURICULAR CANAL|MERKEL CELL CARCINOMA OF LEFT EAR AND EXTERNAL AURIC CANAL
C2857293|T037|S72.123C|ICD10CM|DISPLACED FRACTURE OF LESSER TROCHANTER OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF LESS TROCHANTER OF UNSP FEMR, 7THC
C2857292|T037|S72.123B|ICD10CM|DISPLACED FRACTURE OF LESSER TROCHANTER OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF LESS TROCHANTER OF UNSP FEMR, 7THB
C0031036|T047|M30.0|DMDICD10|POLYARTERITIS NODOSA|PANARTERIITIS NODOSA
C0008728|T047|M30.1|DMDICD10|POLYARTERITIS WITH LUNG INVOLVEMENT [CHURG-STRAUSS]|PANARTERIITIS MIT LUNGENBETEILIGUNG
C0348857|T047|M30.2|DMDICD10|JUVENILE POLYARTERITIS|JUVENILE PANARTERIITIS
C0026691|T047|M30.3|DMDICD10|MUCOCUTANEOUS LYMPH NODE SYNDROME [KAWASAKI]|MUKOKUTANES LYMPHKNOTENSYNDROM [KAWASAKI-KRANKHEIT]
C2838487|T037|S32.699B|ICD10CM|OTHER SPECIFIED FRACTURE OF UNSPECIFIED ISCHIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF UNSP ISCHIUM, INIT ENCNTR FOR OPEN FRACTURE
C0477584|T047|M30.8|DMDICD10|OTHER CONDITIONS RELATED TO POLYARTERITIS NODOSA|SONSTIGE MIT PANARTERIITIS NODOSA VERWANDTE ZUSTAENDE
C2876645|T037|T36.4X2S|ICD10CM|POISONING BY TETRACYCLINES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY TETRACYCLINES, INTENTIONAL SELF-HARM, SEQUELA
C2838179|T037|S32.451A|ICD10CM|DISPLACED TRANSVERSE FRACTURE OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED TRANSVERSE FRACTURE OF RIGHT ACETABULUM, INIT
C2838180|T037|S32.451B|ICD10CM|DISPLACED TRANSVERSE FRACTURE OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISPLACED TRANSVERSE FX RIGHT ACETABULUM, INIT FOR OPN FX
C3264211|T047|H40.1310|ICD10CM|PIGMENTARY GLAUCOMA, RIGHT EYE, STAGE UNSPECIFIED|PIGMENTARY GLAUCOMA, RIGHT EYE, STAGE UNSPECIFIED
C2889285|T047|M05.559|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP|RHEUMATOID POLYNEUROPATHY W RHEUMATOID ARTHRITIS OF UNSP HIP
C3264041|T047|G43.C0|ICD10CM|PERIODIC HEADACHE SYNDROMES IN CHILD OR ADULT, NOT INTRACTABLE|PERIODIC HEADACHE SYNDROMES IN CHILD OR ADULT, WITHOUT REFRACTORY MIGRAINE
C3264042|T047|G43.C1|ICD10CM|PERIODIC HEADACHE SYNDROMES IN CHILD OR ADULT, INTRACTABLE|PERIODIC HEADACHE SYNDROMES IN CHILD OR ADULT, WITH REFRACTORY MIGRAINE
C2885611|T037|T63.412S|ICD10CM|TOXIC EFFECT OF VENOM OF CENTIPEDES AND VENOMOUS MILLIPEDES, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF VENOM OF CENTIPEDE/MILLIPEDE, SLF-HRM, SQLA
C2848419|T037|S58.112A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN ELBOW AND WRIST, LEFT ARM, INITIAL ENCOUNTER|COMPLETE TRAUM AMP AT LEV BETW ELBOW AND WRS, LEFT ARM, INIT
C2855976|T037|S68.511S|ICD10CM|COMPLETE TRAUMATIC TRANSPHALANGEAL AMPUTATION OF RIGHT THUMB, SEQUELA|COMPLETE TRAUMATIC TRNSPHAL AMPUTATION OF R THM, SEQUELA
C2890530|T037|T84.060A|ICD10CM|WEAR OF ARTICULAR BEARING SURFACE OF INTERNAL PROSTHETIC RIGHT HIP JOINT, INITIAL ENCOUNTER|WEAR OF ARTIC BEARING SURFACE OF INT PROSTH R HIP JT, INIT
C2858748|T037|S72.451A|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPL SUPRCNDL FX W/O INTRCNDL EXTN LOWER END R FEMUR, INIT
C2842077|T191|C50.011|ICD10CM|MALIGNANT NEOPLASM OF NIPPLE AND AREOLA, RIGHT FEMALE BREAST|MALIGNANT NEOPLASM OF NIPPLE AND AREOLA, RIGHT FEMALE BREAST
C2858750|T037|S72.451C|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL SUPRCNDL FX W/O INTRCNDL EXTN LOW END R FEMR, 7THC
C2858749|T037|S72.451B|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL SUPRCNDL FX W/O INTRCNDL EXTN LOW END R FEMR, 7THB
C2874111|T047|E11.618|ICD10CM|TYPE 2 DIABETES MELLITUS WITH OTHER DIABETIC ARTHROPATHY|TYPE 2 DIABETES MELLITUS WITH OTHER DIABETIC ARTHROPATHY
C2869897|T037|S98.919S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED FOOT, LEVEL UNSPECIFIED, SEQUELA|COMPLETE TRAUMATIC AMP OF UNSP FOOT, LEVEL UNSP, SEQUELA
C2874110|T047|E11.610|ICD10CM|TYPE 2 DIABETES MELLITUS WITH DIABETIC NEUROPATHIC ARTHROPATHY|TYPE 2 DIABETES MELLITUS W DIABETIC NEUROPATHIC ARTHROPATHY
C2896728|T046|M80.841A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, RIGHT HAND, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, RIGHT HAND, INIT
C2869895|T037|S98.919A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED FOOT, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF UNSP FOOT, LEVEL UNSP, INIT
C2869896|T037|S98.919D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF UNSPECIFIED FOOT, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF UNSP FOOT, LEVEL UNSP, SUBS
C0025268|T191|E31.22|ICD10CM|MULTIPLE ENDOCRINE NEOPLASIA [MEN] TYPE IIA|MULTIPLE ENDOCRINE NEOPLASIA [MEN] TYPE IIA
C2879797|T037|T47.5X2A|ICD10CM|POISONING BY DIGESTANTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY DIGESTANTS, INTENTIONAL SELF-HARM, INIT ENCNTR
C0260763|T033|Z43.3|DMDICD10|ENCOUNTER FOR ATTENTION TO COLOSTOMY|VERSORGUNG EINES KOLOSTOMAS
C2853845|T191|C82.57|ICD10CM|DIFFUSE FOLLICLE CENTER LYMPHOMA, SPLEEN|DIFFUSE FOLLICLE CENTER LYMPHOMA, SPLEEN
C0260761|T033|Z43.1|DMDICD10|ENCOUNTER FOR ATTENTION TO GASTROSTOMY|VERSORGUNG EINES GASTROSTOMAS
C0260760|T033|Z43.0|DMDICD10|ENCOUNTER FOR ATTENTION TO TRACHEOSTOMY|VERSORGUNG EINES TRACHEOSTOMAS
C2910816|T033|Z43.6|ICD10CM|ENCOUNTER FOR ATTENTION TO OTHER ARTIFICIAL OPENINGS OF URINARY TRACT|ENCOUNTER FOR ATTENTION TO URETHROSTOMY
C0260765|T033|Z43.5|DMDICD10|ENCOUNTER FOR ATTENTION TO CYSTOSTOMY|VERSORGUNG EINES ZYSTOSTOMAS
C2854037|T191|C85.24|ICD10CM|MEDIASTINAL (THYMIC) LARGE B-CELL LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB|MEDIASTNL LARGE B-CELL LYMPH, NODES OF AXILLA AND UPPER LIMB
C2883986|T037|T51.0X2A|ICD10CM|TOXIC EFFECT OF ETHANOL, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF ETHANOL, INTENTIONAL SELF-HARM, INIT ENCNTR
C2910819|T033|Z43.8|ICD10CM|ENCOUNTER FOR ATTENTION TO OTHER ARTIFICIAL OPENINGS|ENCOUNTER FOR ATTENTION TO OTHER ARTIFICIAL OPENINGS
C2853843|T191|C82.55|ICD10CM|DIFFUSE FOLLICLE CENTER LYMPHOMA, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|DIFFUS FOLICL CNTR LYMPH, NODES OF ING REGION AND LOWER LIMB
C2848410|T037|S58.029A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT ELBOW LEVEL, UNSPECIFIED ARM, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION AT ELBOW LEVEL, UNSP ARM, INIT
C2853842|T191|C82.54|ICD10CM|DIFFUSE FOLLICLE CENTER LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB|DIFFUSE FOLICL CENTER LYMPH, NODES OF AXILLA AND UPPER LIMB
C2883988|T037|T51.0X2S|ICD10CM|TOXIC EFFECT OF ETHANOL, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF ETHANOL, INTENTIONAL SELF-HARM, SEQUELA
C2853841|T191|C82.53|ICD10CM|DIFFUSE FOLLICLE CENTER LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES|DIFFUSE FOLLICLE CENTER LYMPHOMA, INTRA-ABD LYMPH NODES
C2848412|T037|S58.029S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT ELBOW LEVEL, UNSPECIFIED ARM, SEQUELA|PARTIAL TRAUMATIC AMP AT ELBOW LEVEL, UNSP ARM, SEQUELA
C2854033|T191|C85.20|ICD10CM|MEDIASTINAL (THYMIC) LARGE B-CELL LYMPHOMA, UNSPECIFIED SITE|MEDIASTINAL (THYMIC) LARGE B-CELL LYMPHOMA, UNSPECIFIED SITE
C2884883|T037|T59.3X2S|ICD10CM|TOXIC EFFECT OF LACRIMOGENIC GAS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF LACRIMOGENIC GAS, SELF-HARM, SEQUELA
C2888302|T047|L89.124|ICD10CM|PRESSURE ULCER OF LEFT UPPER BACK, STAGE 4|PRESSURE ULCER OF LEFT UPPER BACK, STAGE 4
C2888296|T047|L89.122|ICD10CM|PRESSURE ULCER OF LEFT UPPER BACK, STAGE 2|PRESSURE ULCER OF LEFT UPPER BACK, STAGE 2
C2888299|T047|L89.123|ICD10CM|PRESSURE ULCER OF LEFT UPPER BACK, STAGE 3|PRESSURE ULCER OF LEFT UPPER BACK, STAGE 3
C2888290|T047||ICD10CM|PRESSURE ULCER OF LEFT UPPER BACK, UNSTAGEABLE
C2888293|T047|L89.121|ICD10CM|PRESSURE ULCER OF LEFT UPPER BACK, STAGE 1|PRESSURE ULCER OF LEFT UPPER BACK, STAGE 1
C4268161|T047|E13.3533|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, BILATERAL|OTH DIAB WITH PROLIF DIAB RTNOP WITH TRCTN DTCH N-MCLA, BI
C4268160|T047|E13.3532|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, LEFT EYE|OTH DIAB W PROLIF DIAB RTNOP WITH TRCTN DTCH N-MCLA, L EYE
C4268159|T047|E13.3531|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH TRACTION RETINAL DETACHMENT NOT INVOLVING THE MACULA, RIGHT EYE|OTH DIAB W PROLIF DIAB RTNOP WITH TRCTN DTCH N-MCLA, R EYE
C2853838|T191|C82.50|ICD10CM|DIFFUSE FOLLICLE CENTER LYMPHOMA, UNSPECIFIED SITE|DIFFUSE FOLLICLE CENTER LYMPHOMA, UNSPECIFIED SITE
C2888305|T047|L89.129|ICD10CM|PRESSURE ULCER OF LEFT UPPER BACK, UNSPECIFIED STAGE|PRESSURE ULCER OF LEFT UPPER BACK, UNSPECIFIED STAGE
C2884881|T037|T59.3X2A|ICD10CM|TOXIC EFFECT OF LACRIMOGENIC GAS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF LACRIMOGENIC GAS, SELF-HARM, INIT
C3263954|T048|F78|ICD10CM|OTHER INTELLECTUAL DISABILITIES|OTHER INTELLECTUAL DISABILITIES
C3161331|T048|F79|ICD10CM|UNSPECIFIED INTELLECTUAL DISABILITIES|UNSPECIFIED INTELLECTUAL DISABILITIES
C2837971|T191|C40.11|ICD10CM|MALIGNANT NEOPLASM OF SHORT BONES OF RIGHT UPPER LIMB|MALIGNANT NEOPLASM OF SHORT BONES OF RIGHT UPPER LIMB
C2837970|T191|C40.10|ICD10CM|MALIGNANT NEOPLASM OF SHORT BONES OF UNSPECIFIED UPPER LIMB|MALIGNANT NEOPLASM OF SHORT BONES OF UNSPECIFIED UPPER LIMB
C2837972|T191|C40.12|ICD10CM|MALIGNANT NEOPLASM OF SHORT BONES OF LEFT UPPER LIMB|MALIGNANT NEOPLASM OF SHORT BONES OF LEFT UPPER LIMB
C2874985|T048|F70|ICD10CM|MILD INTELLECTUAL DISABILITIES|IQ LEVEL 50-55 TO APPROXIMATELY 70
C2874986|T048|F71|ICD10CM|MODERATE INTELLECTUAL DISABILITIES|IQ LEVEL 35-40 TO 50-55
C2874987|T048|F72|ICD10CM|SEVERE INTELLECTUAL DISABILITIES|IQ 20-25 TO 35-40
C3161330|T048|F73|ICD10CM|PROFOUND INTELLECTUAL DISABILITIES|PROFOUND INTELLECTUAL DISABILITIES
C2882876|T047|I70.529|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, UNSPECIFIED EXTREMITY|ATHSCL NONAUT BIO BYPASS OF EXTRM W REST PAIN, UNSP EXTRM
C2882875|T047|I70.528|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, OTHER EXTREMITY|ATHSCL NONAUT BIO BYPASS OF THE EXTRM W REST PAIN, OTH EXTRM
C2882872|T047|I70.521|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, RIGHT LEG|ATHSCL NONAUT BIO BYPASS OF THE EXTRM W REST PAIN, RIGHT LEG
C0340648|T047||ICD10CM|CORONARY ARTERY DISSECTION
C2882171|T020|I25.41|ICD10CM|CORONARY ARTERY ANEURYSM|CORONARY ARTERIOVENOUS FISTULA, ACQUIRED
C2882873|T047|I70.522|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH REST PAIN, LEFT LEG|ATHSCL NONAUT BIO BYPASS OF THE EXTRM W REST PAIN, LEFT LEG
C4270334|T046|T83.591A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO IMPLANTED URINARY SPHINCTER, INITIAL ENCOUNTER|I/I REACT D/T IMPLANTED URINARY SPHINCTER, INITIAL ENCOUNTER
C2869755|T037|S98.011A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT FOOT AT ANKLE LEVEL, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMP OF RIGHT FOOT AT ANKLE LEVEL, INIT
C0032533|T047|M35.3|DMDICD10|POLYMYALGIA RHEUMATICA|POLYMYALGIA RHEUMATICA
C2876195|T037|T32.44|ICD10CM|CORROSIONS INVOLVING 40-49% OF BODY SURFACE WITH 40-49% THIRD DEGREE CORROSION|CORROS 40-49% OF BODY SURFACE W 40-49% THIRD DEGREE CORROS
C2833876|T037|S14.108S|ICD10CM|UNSPECIFIED INJURY AT C8 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|UNSP INJURY AT C8 LEVEL OF CERVICAL SPINAL CORD, SEQUELA
C2876193|T037|T32.42|ICD10CM|CORROSIONS INVOLVING 40-49% OF BODY SURFACE WITH 20-29% THIRD DEGREE CORROSION|CORROS 40-49% OF BODY SURFACE W 20-29% THIRD DEGREE CORROS
C2902434|T047|M90.532|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, LEFT FOREARM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, LEFT FOREARM
C2832604|T037|S06.823S|ICD10CM|INJURY OF LEFT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, SEQUELA|INJ L INT CAROTID, INTCR W LOC OF 1-5 HRS 59 MIN, SEQUELA
C2832194|T037|S06.334A|ICD10CM|CONTUSION AND LACERATION OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|CONTUS/LAC CEREB, W LOC OF 6 HOURS TO 24 HOURS, INIT
C0477590|T047|M35.1|DMDICD10|OTHER OVERLAP SYNDROMES|SONSTIGE OVERLAP-SYNDROME
C0348257|T047|B39.2|DMDICD10|PULMONARY HISTOPLASMOSIS CAPSULATI, UNSPECIFIED|HISTOPLASMOSE DER LUNGE DURCH HISTOPLASMA CAPSULATUM, NICHT NAEHER BEZEICHNET
C2869757|T037|S98.011S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF RIGHT FOOT AT ANKLE LEVEL, SEQUELA|COMPLETE TRAUMATIC AMP OF RIGHT FOOT AT ANKLE LEVEL, SEQUELA
C2832602|T037|S06.823A|ICD10CM|INJURY OF LEFT INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION, NOT ELSEWHERE CLASSIFIED WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|INJURY OF L INT CAROTID, INTCR W LOC OF 1-5 HRS 59 MIN, INIT
C4269256|T037|S02.110S|ICD10CM|TYPE I OCCIPITAL CONDYLE FRACTURE, UNSPECIFIED SIDE, SEQUELA|TYPE I OCCIPITAL CONDYLE FRACTURE, UNSPECIFIED SIDE, SEQUELA
C0343899|T047|B39.1|DMDICD10|CHRONIC PULMONARY HISTOPLASMOSIS CAPSULATI|CHRONISCHE HISTOPLASMOSE DER LUNGE DURCH HISTOPLASMA CAPSULATUM
C4269251|T037|S02.110A|ICD10CM|TYPE I OCCIPITAL CONDYLE FRACTURE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE I OCCIPITAL CONDYLE FRACTURE, UNSPECIFIED SIDE, INIT
C4269252|T037|S02.110B|ICD10CM|TYPE I OCCIPITAL CONDYLE FRACTURE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE I OCCIPITAL CONDYLE FRACTURE, UNSPECIFIED SIDE, 7THB
C2902435|T047|M90.539|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, UNSPECIFIED FOREARM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, UNSP FOREARM
C2835392|T037|S22.068B|ICD10CM|OTHER FRACTURE OF T7-T8 THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF T7-T8 THORACIC VERTEBRA, INIT FOR OPN FX
C2835391|T037|S22.068A|ICD10CM|OTHER FRACTURE OF T7-T8 THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF T7-T8 THORACIC VERTEBRA, INIT FOR CLOS FX
C2833272|T037|S12.131B|ICD10CM|UNSPECIFIED TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP TRAUM NONDISP SPONDYLOLYSIS OF 2ND CERVCAL VERT, 7THB
C2901783|T047|M86.051|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, RIGHT FEMUR|ACUTE HEMATOGENOUS OSTEOMYELITIS, RIGHT FEMUR
C2901784|T047|M86.052|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, LEFT FEMUR|ACUTE HEMATOGENOUS OSTEOMYELITIS, LEFT FEMUR
C2833271|T037|S12.131A|ICD10CM|UNSPECIFIED TRAUMATIC NONDISPLACED SPONDYLOLISTHESIS OF SECOND CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP TRAUM NONDISP SPONDYLOLYSIS OF 2ND CERVCAL VERT, INIT
C2905663|T037|X71.8XXD|ICD10CM|OTHER INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION, SUBSEQUENT ENCOUNTER|OTH INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION, SUBS
C2901785|T047|M86.059|ICD10CM|ACUTE HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED FEMUR|ACUTE HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED FEMUR
C2874841|T048|F19.930|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH WITHDRAWAL, UNCOMPLICATED|OTH PSYCHOACTIVE SUBSTANCE USE, UNSP W WITHDRAWAL, UNCOMP
C2889477|T047|M06.839|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, UNSPECIFIED WRIST|OTHER SPECIFIED RHEUMATOID ARTHRITIS, UNSPECIFIED WRIST
C2848447|T037|S58.912S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT FOREARM, LEVEL UNSPECIFIED, SEQUELA|COMPLETE TRAUMATIC AMP OF L FOREARM, LEVEL UNSP, SEQUELA
C2843305|T037|S48.119S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN UNSPECIFIED SHOULDER AND ELBOW, SEQUELA|COMPLETE TRAUM AMP AT LEVEL BETW UNSP SHLDR AND ELBOW, SQLA
C2885784|T037|T63.622S|ICD10CM|TOXIC EFFECT OF CONTACT WITH OTHER JELLYFISH, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CONTACT W OTH JELLYFISH, SELF-HARM, SEQUELA
C2905812|T037|X83.1XXS|ICD10CM|INTENTIONAL SELF-HARM BY ELECTROCUTION, SEQUELA|INTENTIONAL SELF-HARM BY ELECTROCUTION, SEQUELA
C2885782|T037|T63.622A|ICD10CM|TOXIC EFFECT OF CONTACT WITH OTHER JELLYFISH, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CONTACT W OTH JELLYFISH, SELF-HARM, INIT
C2848445|T037|S58.912A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT FOREARM, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF L FOREARM, LEVEL UNSP, INIT
C2889617|T047|M08.859|ICD10CM|OTHER JUVENILE ARTHRITIS, UNSPECIFIED HIP|OTHER JUVENILE ARTHRITIS, UNSPECIFIED HIP
C2905811|T037|X83.1XXD|ICD10CM|INTENTIONAL SELF-HARM BY ELECTROCUTION, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY ELECTROCUTION, SUBSEQUENT ENCOUNTER
C2889616|T047|M08.852|ICD10CM|OTHER JUVENILE ARTHRITIS, LEFT HIP|OTHER JUVENILE ARTHRITIS, LEFT HIP
C2905810|T037|X83.1XXA|ICD10CM|INTENTIONAL SELF-HARM BY ELECTROCUTION, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY ELECTROCUTION, INITIAL ENCOUNTER
C2889615|T047|M08.851|ICD10CM|OTHER JUVENILE ARTHRITIS, RIGHT HIP|OTHER JUVENILE ARTHRITIS, RIGHT HIP
C0348989|T047|B44.2|DMDICD10|TONSILLAR ASPERGILLOSIS|ASPERGILLOSE DER TONSILLEN
C2501343|T060|B440|ICD10PCS|INVASIVE PULMONARY ASPERGILLOSIS|IMAGING @ LOWER ARTERIES @ ULTRASONOGRAPHY @ ABDOMINAL AORTA
C0348258|T047|B44.1|DMDICD10|OTHER PULMONARY ASPERGILLOSIS|SONSTIGE ASPERGILLOSE DER LUNGE
C2501355|T060|B447|ICD10PCS|DISSEMINATED ASPERGILLOSIS|IMAGING @ LOWER ARTERIES @ ULTRASONOGRAPHY @ RENAL ARTERY, LEFT
C2833488|T037|S12.450B|ICD10CM|OTHER TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF FIFTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH TRAUM DISPL SPONDYLOLYSIS OF 5TH CERVCAL VERT, 7THB
C0004030|T047|B44.9|DMDICD10|ASPERGILLOSIS, UNSPECIFIED|ASPERGILLOSE, NICHT NAEHER BEZEICHNET
C2889223|T047|M05.369|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP KNEE
C2889360|T047|M05.819|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED SHOULDER|OTH RHEU ARTHRITIS W RHEUMATOID FACTOR OF UNSP SHOULDER
C2889222|T047|M05.362|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT KNEE|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889221|T047|M05.361|ICD10CM|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT KNEE|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889358|T047|M05.811|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT SHOULDER|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF R SHOULDER
C2832647|T037|S06.894A|ICD10CM|OTHER SPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS, INITIAL ENCOUNTER|INTCRAN INJ W LOC OF 6 HOURS TO 24 HOURS, INIT
C2889359|T047|M05.812|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT SHOULDER|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF L SHOULDER
C2887137|T047|I82.A11|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF RIGHT AXILLARY VEIN|ACUTE EMBOLISM AND THROMBOSIS OF RIGHT AXILLARY VEIN
C2887139|T047|I82.A13|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF AXILLARY VEIN, BILATERAL|ACUTE EMBOLISM AND THROMBOSIS OF AXILLARY VEIN, BILATERAL
C2887138|T047|I82.A12|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF LEFT AXILLARY VEIN|ACUTE EMBOLISM AND THROMBOSIS OF LEFT AXILLARY VEIN
C2887140|T047|I82.A19|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED AXILLARY VEIN|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED AXILLARY VEIN
C2874813|T048|F19.221|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH INTOXICATION DELIRIUM|OTH PSYCHOACTIVE SUBSTANCE DEPENDENCE W INTOX DELIRIUM
C0348636|T046|I63.8|DMDICD10|OTHER CEREBRAL INFARCTION|SONSTIGER HIRNINFARKT
C0038454|T047||ICD10CM|CEREBRAL INFARCTION, UNSPECIFIED
C2833964|T037|S14.133A|ICD10CM|ANTERIOR CORD SYNDROME AT C3 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|ANTERIOR CORD SYNDROME AT C3, INIT
C2859156|T037|S73.005A|ICD10CM|UNSPECIFIED DISLOCATION OF LEFT HIP, INITIAL ENCOUNTER|UNSPECIFIED DISLOCATION OF LEFT HIP, INITIAL ENCOUNTER
C2855919|T037|S68.123S|ICD10CM|PARTIAL TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF LEFT MIDDLE FINGER, SEQUELA|PARTIAL TRAUMATIC MCP AMPUTATION OF L MID FINGER, SEQUELA
C2833965|T037|S14.133D|ICD10CM|ANTERIOR CORD SYNDROME AT C3 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|ANTERIOR CORD SYNDROME AT C3, SUBS
C2832325|T037|S06.365A|ICD10CM|TRAUMATIC HEMORRHAGE OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, INITIAL ENCOUNTER|TRAUM HEMOR CEREB, W LOC >24 HR W RET CONSC LEV, INIT
C0451676|T047|I63.6|DMDICD10|CEREBRAL INFARCTION DUE TO CEREBRAL VENOUS THROMBOSIS, NONPYOGENIC|HIRNINFARKT DURCH THROMBOSE DER HIRNVENEN, NICHTEITRIG
C2833966|T037|S14.133S|ICD10CM|ANTERIOR CORD SYNDROME AT C3 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|ANTERIOR CORD SYNDROME AT C3, SEQUELA
C2838272|T037|S32.472A|ICD10CM|DISPLACED FRACTURE OF MEDIAL WALL OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF MEDIAL WALL OF LEFT ACETABULUM, INIT FOR CLOS FX
C2833929|T037|S14.123S|ICD10CM|CENTRAL CORD SYNDROME AT C3 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|CENTRAL CORD SYNDROME AT C3, SEQUELA
C2878121|T037|T42.3X2A|ICD10CM|POISONING BY BARBITURATES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY BARBITURATES, INTENTIONAL SELF-HARM, INIT
C2883088|T047|I82.290|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF OTHER THORACIC VEINS|ACUTE EMBOLISM AND THROMBOSIS OF OTHER THORACIC VEINS
C2883089|T047|I82.291|ICD10CM|CHRONIC EMBOLISM AND THROMBOSIS OF OTHER THORACIC VEINS|CHRONIC EMBOLISM AND THROMBOSIS OF OTHER THORACIC VEINS
C2877382|T037|T39.1X2A|ICD10CM|POISONING BY 4-AMINOPHENOL DERIVATIVES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY 4-AMINOPHENOL DERIVATIVES, SELF-HARM, INIT
C2869867|T037|S98.312S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT MIDFOOT, SEQUELA|COMPLETE TRAUMATIC AMPUTATION OF LEFT MIDFOOT, SEQUELA
C2884334|T037|T53.92XA|ICD10CM|TOXIC EFFECT OF UNSPECIFIED HALOGEN DERIVATIVES OF ALIPHATIC AND AROMATIC HYDROCARBONS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOX EFF OF UNSP HALGN DERIV OF AROMAT HYDROCRB,SLF-HRM, INIT
C2890111|T037|T82.593A|ICD10CM|OTHER MECHANICAL COMPLICATION OF BALLOON (COUNTERPULSATION) DEVICE, INITIAL ENCOUNTER|MECH COMPL OF BALLOON (COUNTERPULSATION) DEVICE, INIT ENCNTR
C2869865|T037|S98.312A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT MIDFOOT, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF LEFT MIDFOOT, INIT ENCNTR
C2887488|T047|J86.9|ICD10CM|PYOTHORAX WITHOUT FISTULA|EMPYEMA (CHEST) (LUNG) (PLEURA)
C2869866|T037|S98.312D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT MIDFOOT, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF LEFT MIDFOOT, SUBS ENCNTR
C2887487|T047|J86.0|ICD10CM|PYOTHORAX WITH FISTULA|ANY CONDITION CLASSIFIABLE TO J86.9 WITH FISTULA
C2885765|T037|T63.612A|ICD10CM|TOXIC EFFECT OF CONTACT WITH PORTUGESE MAN-O-WAR, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF CONTACT W PORTUGESE MAN-O-WAR, SLF-HRM, INIT
C2832327|T037|S06.365S|ICD10CM|TRAUMATIC HEMORRHAGE OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, SEQUELA|TRAUM HEMOR CEREB, W LOC >24 HR W RET CONSC LEV, SEQUELA
C0154683|T047|G12.29|ICD10CM|OTHER MOTOR NEURON DISEASE|OTHER MOTOR NEURON DISEASE
C4082951|T047|G12.25|ICD10CM|PROGRESSIVE SPINAL MUSCLE ATROPHY|PROGRESSIVE SPINAL MUSCLE ATROPHY
C0270763|T047||ICD10CM|FAMILIAL MOTOR NEURON DISEASE
C0002736|T047||ICD10CM|AMYOTROPHIC LATERAL SCLEROSIS
C0085084|T047|G12.20|ICD10CM|MOTOR NEURON DISEASE, UNSPECIFIED|MOTOR NEURON DISEASE, UNSPECIFIED
C0154682|T047||ICD10CM|PRIMARY LATERAL SCLEROSIS
C0030442|T047|G12.22|ICD10CM|PROGRESSIVE BULBAR PALSY|PROGRESSIVE BULBAR PALSY
C1510446|T047|I24.9|DMDICD10|ACUTE ISCHEMIC HEART DISEASE, UNSPECIFIED|AKUTE ISCHAEMISCHE HERZKRANKHEIT, NICHT NAEHER BEZEICHNET
C0348590|T047|I24|DMDICD10|OTHER FORMS OF ACUTE ISCHEMIC HEART DISEASE|SONSTIGE AKUTE ISCHAEMISCHE HERZKRANKHEIT
C4236949|T048|F10.959|ICD10CM|ALCOHOL USE, UNSPECIFIED WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|ALCOHOL-INDUCED PSYCHOTIC DISORDER WITHOUT USE DISORDER
C2878123|T037|T42.3X2S|ICD10CM|POISONING BY BARBITURATES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY BARBITURATES, INTENTIONAL SELF-HARM, SEQUELA
C0152107|T047|I24.1|DMDICD10|DRESSLER'S SYNDROME|POSTMYOKARDINFARKT-SYNDROM
C2882160|T047|I24.0|ICD10CM|ACUTE CORONARY THROMBOSIS NOT RESULTING IN MYOCARDIAL INFARCTION|ACUTE CORONARY THROMBOSIS NOT RESULTING IN MYOCARDIAL INFRC
C2874412|T048|F10.951|ICD10CM|ALCOHOL USE, UNSPECIFIED WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|ALCOHOL USE, UNSP W ALCOH-INDUCE PSYCH DISORDER W HALLUCIN
C2874411|T048|F10.950|ICD10CM|ALCOHOL USE, UNSPECIFIED WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|ALCOHOL USE, UNSP W ALCOH-INDUCE PSYCH DISORDER W DELUSIONS
C2869884|T037|S98.329S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED MIDFOOT, SEQUELA|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED MIDFOOT, SEQUELA
C2884996|T037|T59.92XS|ICD10CM|TOXIC EFFECT OF UNSPECIFIED GASES, FUMES AND VAPORS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF UNSP GASES, FUMES AND VAPORS, SLF-HRM, SQLA
C2901068|T046|M84.472A|ICD10CM|PATHOLOGICAL FRACTURE, LEFT ANKLE, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, LEFT ANKLE, INIT ENCNTR FOR FRACTURE
C2869883|T037|S98.329D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED MIDFOOT, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF UNSP MIDFOOT, SUBS ENCNTR
C2869882|T037|S98.329A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED MIDFOOT, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF UNSP MIDFOOT, INIT ENCNTR
C0153491|T191|C34.2|DMDICD10|MALIGNANT NEOPLASM OF MIDDLE LOBE, BRONCHUS OR LUNG|BOESARTIGE NEUBILDUNG: MITTELLAPPEN (-BRONCHUS)
C2884994|T037|T59.92XA|ICD10CM|TOXIC EFFECT OF UNSPECIFIED GASES, FUMES AND VAPORS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF UNSP GASES, FUMES AND VAPORS, SLF-HRM, INIT
C2874122|T047||ICD10CM|TYPE 2 DIABETES MELLITUS WITH HYPOGLYCEMIA WITHOUT COMA
C2902371|T047|M89.649|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, UNSPECIFIED HAND|OSTEOPATHY AFTER POLIOMYELITIS, UNSPECIFIED HAND
C2889400|T047|M06.049|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, UNSPECIFIED HAND|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, UNSP HAND
C2889399|T047|M06.042|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, LEFT HAND|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, LEFT HAND
C2889398|T047|M06.041|ICD10CM|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, RIGHT HAND|RHEUMATOID ARTHRITIS WITHOUT RHEUMATOID FACTOR, RIGHT HAND
C4509243|T047|I50.814|ICD10CM|RIGHT HEART FAILURE DUE TO LEFT HEART FAILURE|RIGHT VENTRICULAR FAILURE SECONDARY TO LEFT VENTRICULAR FAILURE
C4509241|T047|I50.813|ICD10CM|ACUTE ON CHRONIC RIGHT HEART FAILURE|ACUTE EXACERBATION OF CHRONIC (ISOLATED) RIGHT VENTRICULAR FAILURE
C4509236|T047|I50.812|ICD10CM|CHRONIC RIGHT HEART FAILURE|CHRONIC (ISOLATED) RIGHT VENTRICULAR FAILURE
C4509233|T047|I50.811|ICD10CM|ACUTE RIGHT HEART FAILURE|ACUTE (ISOLATED) RIGHT VENTRICULAR FAILURE
C4509231|T047|I50.810|ICD10CM|RIGHT HEART FAILURE, UNSPECIFIED|RIGHT HEART FAILURE WITHOUT MENTION OF LEFT HEART FAILURE
C0451670|T047|G70.2|DMDICD10|CONGENITAL AND DEVELOPMENTAL MYASTHENIA|ANGEBORENE ODER ENTWICKLUNGSBEDINGTE MYASTHENIE
C2834010|T037|S14.145D|ICD10CM|BROWN-SEQUARD SYNDROME AT C5 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|BROWN-SEQUARD SYNDROME AT C5, SUBS
C4269473|T037|S02.621S|ICD10CM|FRACTURE OF SUBCONDYLAR PROCESS OF RIGHT MANDIBLE, SEQUELA|FRACTURE OF SUBCONDYLAR PROCESS OF RIGHT MANDIBLE, SEQUELA
C2875137|T047|G40.89|ICD10CM|OTHER SEIZURES|OTHER SEIZURES
C0393939|T047|G70.1|DMDICD10|TOXIC MYONEURAL DISORDERS|TOXISCHE NEUROMUSKULAERE KRANKHEITEN
C2905775|T037|X80.XXXS|ICD10CM|INTENTIONAL SELF-HARM BY JUMPING FROM A HIGH PLACE, SEQUELA|INTENTIONAL SELF-HARM BY JUMPING FROM A HIGH PLACE, SEQUELA
C2833933|T037|S14.124S|ICD10CM|CENTRAL CORD SYNDROME AT C4 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|CENTRAL CORD SYNDROME AT C4, SEQUELA
C2832103|T037|S06.312A|ICD10CM|CONTUSION AND LACERATION OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|CONTUS/LAC RIGHT CEREBRUM W LOC OF 31-59 MIN, INIT
C2905774|T037|X80.XXXD|ICD10CM|INTENTIONAL SELF-HARM BY JUMPING FROM A HIGH PLACE, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY JUMPING FROM A HIGH PLACE, SUBS
C2835263|T037|S22.030B|ICD10CM|WEDGE COMPRESSION FRACTURE OF THIRD THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|WEDGE COMPRSN FX THIRD THOR VERTEBRA, INIT FOR OPN FX
C2835262|T037|S22.030A|ICD10CM|WEDGE COMPRESSION FRACTURE OF THIRD THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|WEDGE COMPRESSION FRACTURE OF THIRD THORACIC VERTEBRA, INIT
C0349080|T048|G10|ICD10CM|HUNTINGTON'S DISEASE|HUNTINGTON'S DEMENTIA
C4509349|T047|M33.02|ICD10CM|JUVENILE DERMATOMYOSITIS WITH MYOPATHY|JUVENILE DERMATOMYOSITIS WITH MYOPATHY
C4509350|T047|M33.03|ICD10CM|JUVENILE DERMATOMYOSITIS WITHOUT MYOPATHY|JUVENILE DERMATOMYOSITIS WITHOUT MYOPATHY
C4509347|T047|M33.00|ICD10CM|JUVENILE DERMATOMYOSITIS, ORGAN INVOLVEMENT UNSPECIFIED|JUVENILE DERMATOMYOSITIS, ORGAN INVOLVEMENT UNSPECIFIED
C4509348|T047|M33.01|ICD10CM|JUVENILE DERMATOMYOSITIS WITH RESPIRATORY INVOLVEMENT|JUVENILE DERMATOMYOSITIS WITH RESPIRATORY INVOLVEMENT
C2837706|T037|S32.121A|ICD10CM|MINIMALLY DISPLACED ZONE II FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|MINIMALLY DISPLACED ZONE II FRACTURE OF SACRUM, INIT
C2837707|T037|S32.121B|ICD10CM|MINIMALLY DISPLACED ZONE II FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|MINIMALLY DISPLACED ZONE II FX SACRUM, INIT FOR OPN FX
C4509587|T047|M33.09|ICD10CM|JUVENILE DERMATOMYOSITIS WITH OTHER ORGAN INVOLVEMENT|JUVENILE DERMATOMYOSITIS WITH OTHER ORGAN INVOLVEMENT
C2875324|T047|G80.3|ICD10CM|ATHETOID CEREBRAL PALSY|DYSTONIC CEREBRAL PALSY
C2853812|T191|C82.26|ICD10CM|FOLLICULAR LYMPHOMA GRADE III, UNSPECIFIED, INTRAPELVIC LYMPH NODES|FOLLICULAR LYMPHOMA GRADE III, UNSP, INTRAPELVIC LYMPH NODES
C2853813|T191|C82.27|ICD10CM|FOLLICULAR LYMPHOMA GRADE III, UNSPECIFIED, SPLEEN|FOLLICULAR LYMPHOMA GRADE III, UNSPECIFIED, SPLEEN
C2853810|T191|C82.24|ICD10CM|FOLLICULAR LYMPHOMA GRADE III, UNSPECIFIED, LYMPH NODES OF AXILLA AND UPPER LIMB|FOLICLAR LYMPH GRADE III, UNSP, NODES OF AXLA AND UPPER LIMB
C2853811|T191|C82.25|ICD10CM|FOLLICULAR LYMPHOMA GRADE III, UNSPECIFIED, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|FOLICLAR LYMPH GRADE III, UNSP, NODES OF ING RGN AND LOW LMB
C2853808|T191|C82.22|ICD10CM|FOLLICULAR LYMPHOMA GRADE III, UNSPECIFIED, INTRATHORACIC LYMPH NODES|FOLLICULAR LYMPHOMA GRADE III, UNSP, INTRATHORAC LYMPH NODES
C2853809|T191|C82.23|ICD10CM|FOLLICULAR LYMPHOMA GRADE III, UNSPECIFIED, INTRA-ABDOMINAL LYMPH NODES|FOLLICULAR LYMPHOMA GRADE III, UNSP, INTRA-ABD LYMPH NODES
C2853806|T191|C82.20|ICD10CM|FOLLICULAR LYMPHOMA GRADE III, UNSPECIFIED, UNSPECIFIED SITE|FOLLICULAR LYMPHOMA GRADE III, UNSPECIFIED, UNSPECIFIED SITE
C2853807|T191|C82.21|ICD10CM|FOLLICULAR LYMPHOMA GRADE III, UNSPECIFIED, LYMPH NODES OF HEAD, FACE, AND NECK|FOLICLAR LYMPH GRADE III, UNSP, NODES OF HEAD, FACE, AND NK
C2831978|T037|S06.1X1S|ICD10CM|TRAUMATIC CEREBRAL EDEMA WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|TRAUM CEREBRAL EDEMA W LOC OF 30 MINUTES OR LESS, SEQUELA
C2837904|T037|S32.409A|ICD10CM|UNSPECIFIED FRACTURE OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF UNSP ACETABULUM, INIT FOR CLOS FX
C2873886|T047|E08.11|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH KETOACIDOSIS WITH COMA|DIABETES DUE TO UNDERLYING CONDITION W KETOACIDOSIS W COMA
C2873885|T047|E08.10|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH KETOACIDOSIS WITHOUT COMA|DIABETES DUE TO UNDERLYING CONDITION W KETOACIDOSIS W/O COMA
C0477735|T047|N15.8|DMDICD10|OTHER SPECIFIED RENAL TUBULO-INTERSTITIAL DISEASES|SONSTIGE NAEHER BEZEICHNETE TUBULOINTERSTITIELLE NIERENKRANKHEITEN
C2875325|T047|G80.8|ICD10CM|OTHER CEREBRAL PALSY|MIXED CEREBRAL PALSY SYNDROMES
C0004698|T047|N15.0|DMDICD10|BALKAN NEPHROPATHY|BALKAN-NEPHROPATHIE
C2831976|T037|S06.1X1A|ICD10CM|TRAUMATIC CEREBRAL EDEMA WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|TRAUMATIC CEREBRAL EDEMA W LOC OF 30 MINUTES OR LESS, INIT
C0023374|T047|E79.1|DMDICD10|LESCH-NYHAN SYNDROME|LESCH-NYHAN-SYNDROM
C2857173|T037|S72.112C|ICD10CM|DISPLACED FRACTURE OF GREATER TROCHANTER OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF GREATER TROCHANTER OF L FEMR, 7THC
C2857172|T037|S72.112B|ICD10CM|DISPLACED FRACTURE OF GREATER TROCHANTER OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF GREATER TROCHANTER OF L FEMR, 7THB
C2857171|T037|S72.112A|ICD10CM|DISPLACED FRACTURE OF GREATER TROCHANTER OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF GREATER TROCHANTER OF LEFT FEMUR, INIT
C2859206|T037|S73.026A|ICD10CM|OBTURATOR DISLOCATION OF UNSPECIFIED HIP, INITIAL ENCOUNTER|OBTURATOR DISLOCATION OF UNSPECIFIED HIP, INITIAL ENCOUNTER
C2848397|T037|S58.019A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT ELBOW LEVEL, UNSPECIFIED ARM, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION AT ELBOW LEVEL, UNSP ARM, INIT
C3263897|T037|T81.11XA|ICD10CM|POSTPROCEDURAL  CARDIOGENIC SHOCK, INITIAL ENCOUNTER|POSTPROCEDURAL CARDIOGENIC SHOCK, INITIAL ENCOUNTER
C0220988|T047|E79.8|ICD10CM|OTHER DISORDERS OF PURINE AND PYRIMIDINE METABOLISM|HEREDITARY XANTHINURIA
C2848399|T037|S58.019S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT ELBOW LEVEL, UNSPECIFIED ARM, SEQUELA|COMPLETE TRAUMATIC AMP AT ELBOW LEVEL, UNSP ARM, SEQUELA
C0472777|T047||ICD10CM|HEMOGLOBIN E-BETA THALASSEMIA
C2877281|T037|T38.902S|ICD10CM|POISONING BY UNSPECIFIED HORMONE ANTAGONISTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY UNSP HORMONE ANTAGONISTS, SELF-HARM, SEQUELA
C2901836|T047|M86.269|ICD10CM|SUBACUTE OSTEOMYELITIS, UNSPECIFIED TIBIA AND FIBULA|SUBACUTE OSTEOMYELITIS, UNSPECIFIED TIBIA AND FIBULA
C0838532|T047|M46.59|ICD10CM|OTHER INFECTIVE SPONDYLOPATHIES, MULTIPLE SITES IN SPINE|OTHER INFECTIVE SPONDYLOPATHIES, MULTIPLE SITES IN SPINE
C0838540|T047|M46.58|ICD10CM|OTHER INFECTIVE SPONDYLOPATHIES, SACRAL AND SACROCOCCYGEAL REGION|OTH INFECTIVE SPONDYLOPATHIES, SACR/SACROCYGL REGION
C0838537|T047|M46.55|ICD10AM|OTHER INFECTIVE SPONDYLOPATHIES, THORACOLUMBAR REGION|OTHER INFECTIVE SPONDYLOPATHIES, THORACOLUMBAR REGION
C0838536|T047|M46.54|ICD10AM|OTHER INFECTIVE SPONDYLOPATHIES, THORACIC REGION|OTHER INFECTIVE SPONDYLOPATHIES, THORACIC REGION
C0838539|T047|M46.57|ICD10AM|OTHER INFECTIVE SPONDYLOPATHIES, LUMBOSACRAL REGION|OTHER INFECTIVE SPONDYLOPATHIES, LUMBOSACRAL REGION
C0838538|T047|M46.56|ICD10AM|OTHER INFECTIVE SPONDYLOPATHIES, LUMBAR REGION|OTHER INFECTIVE SPONDYLOPATHIES, LUMBAR REGION
C0838533|T047|M46.51|ICD10CM|OTHER INFECTIVE SPONDYLOPATHIES, OCCIPITO-ATLANTO-AXIAL REGION|OTH INFECTIVE SPONDYLOPATHIES, OCCIPITO-ATLANTO-AXIAL REGION
C0838532|T047|M46.50|ICD10AM|OTHER INFECTIVE SPONDYLOPATHIES, SITE UNSPECIFIED|OTHER INFECTIVE SPONDYLOPATHIES, MULTIPLE SITES IN SPINE
C0838535|T047|M46.53|ICD10AM|OTHER INFECTIVE SPONDYLOPATHIES, CERVICOTHORACIC REGION|OTHER INFECTIVE SPONDYLOPATHIES, CERVICOTHORACIC REGION
C0838534|T047|M46.52|ICD10AM|OTHER INFECTIVE SPONDYLOPATHIES, CERVICAL REGION|OTHER INFECTIVE SPONDYLOPATHIES, CERVICAL REGION
C2886768|T037|T79.A29A|ICD10CM|TRAUMATIC COMPARTMENT SYNDROME OF UNSPECIFIED LOWER EXTREMITY, INITIAL ENCOUNTER|TRAUMATIC COMPARTMENT SYNDROME OF UNSP LOWER EXTREMITY, INIT
C3161373|T047||ICD10CM|OTHER THALASSEMIAS
C2874509|T048|F12.99|ICD10CM|CANNABIS USE, UNSPECIFIED WITH UNSPECIFIED CANNABIS-INDUCED DISORDER|CANNABIS USE, UNSP WITH UNSP CANNABIS-INDUCED DISORDER
C2875182|T047|G43.811|ICD10CM|OTHER MIGRAINE, INTRACTABLE, WITH STATUS MIGRAINOSUS|OTHER MIGRAINE, INTRACTABLE, WITH STATUS MIGRAINOSUS
C2873965|T047|E09.311|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH UNSPECIFIED DIABETIC RETINOPATHY WITH MACULAR EDEMA|DRUG/CHEM DIABETES W UNSP DIABETIC RTNOP W MACULAR EDEMA
C2873966|T047|E09.319|ICD10CM|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS WITH UNSPECIFIED DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA|DRUG/CHEM DIABETES W UNSP DIABETIC RTNOP W/O MACULAR EDEMA
C0839968|T047|M86.40|ICD10AM|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, UNSPECIFIED SITE|CHRONIC OSTEOMYELITIS WITH DRAINING SINUS, MULTIPLE SITES
C2889572|T047|M08.28|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, VERTEBRAE|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, VERTEBRAE
C2889573|T047|M08.29|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, MULTIPLE SITES|JUVENILE RHEU ARTHRITIS W SYSTEMIC ONSET, MULTIPLE SITES
C1384600|T047|M08.20|ICD10CM|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, UNSPECIFIED SITE|JUVENILE RHEUMATOID ARTHRITIS WITH SYSTEMIC ONSET, UNSPECIFIED SITE
C2889585|T047|M08.441|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, RIGHT HAND|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, RIGHT HAND
C2889586|T047|M08.442|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, LEFT HAND|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, LEFT HAND
C2833982|T037|S14.137S|ICD10CM|ANTERIOR CORD SYNDROME AT C7 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|ANTERIOR CORD SYNDROME AT C7, SEQUELA
C2889587|T047|M08.449|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED HAND|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, UNSP HAND
C2856078|T037|S68.628S|ICD10CM|PARTIAL TRAUMATIC TRANSPHALANGEAL AMPUTATION OF OTHER FINGER, SEQUELA|PARTIAL TRAUMATIC TRNSPHAL AMPUTATION OF FINGER, SEQUELA
C2833228|T037|S12.110B|ICD10CM|ANTERIOR DISPLACED TYPE II DENS FRACTURE, INITIAL ENCOUNTER FOR OPEN FRACTURE|ANTERIOR DISPLACED TYPE II DENS FRACTURE, INIT FOR OPN FX
C2833227|T037|S12.110A|ICD10CM|ANTERIOR DISPLACED TYPE II DENS FRACTURE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|ANTERIOR DISPLACED TYPE II DENS FRACTURE, INIT FOR CLOS FX
C0477325|T047|D82.8|DMDICD10|IMMUNODEFICIENCY ASSOCIATED WITH OTHER SPECIFIED MAJOR DEFECTS|IMMUNDEFEKTE IN VERBINDUNG MIT ANDEREN NAEHER BEZEICHNETEN SCHWEREN DEFEKTEN
C0477326|T047|D82.9|DMDICD10|IMMUNODEFICIENCY ASSOCIATED WITH MAJOR DEFECT, UNSPECIFIED|IMMUNDEFEKT IN VERBINDUNG MIT SCHWEREM DEFEKT, NICHT NAEHER BEZEICHNET
C3887645|T047|D82.4|DMDICD10|HYPERIMMUNOGLOBULIN E [IGE] SYNDROME|HYPERIMMUNGLOBULIN-E[IGE]-SYNDROM
C0265299|T047|D82.2|DMDICD10|IMMUNODEFICIENCY WITH SHORT-LIMBED STATURE|IMMUNDEFEKT MIT DISPROPORTIONIERTEM MINDERWUCHS
C0549463|T191||ICD10CM|IMMUNODEFICIENCY FOLLOWING HEREDITARY DEFECTIVE RESPONSE TO EPSTEIN-BARR VIRUS
C2531321|T061|D820|ICD10PCS|WISKOTT-ALDRICH SYNDROME|RADIATION THERAPY @ EYE @ STEREOTACTIC RADIOSURGERY @ EYE
C2873847|T047|D82.1|ICD10CM|DI GEORGE'S SYNDROME|THYMIC APLASIA OR HYPOPLASIA WITH IMMUNODEFICIENCY
C2878712|T037|T43.92XA|ICD10CM|POISONING BY UNSPECIFIED PSYCHOTROPIC DRUG, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY UNSP PSYCHOTROPIC DRUG, SELF-HARM, INIT
C2890592|T037|T84.113A|ICD10CM|BREAKDOWN (MECHANICAL) OF INTERNAL FIXATION DEVICE OF BONE OF LEFT FOREARM, INITIAL ENCOUNTER|BREAKDOWN OF INT FIX OF BONE OF LEFT FOREARM, INIT
C2878714|T037|T43.92XS|ICD10CM|POISONING BY UNSPECIFIED PSYCHOTROPIC DRUG, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY UNSP PSYCHOTROPIC DRUG, SELF-HARM, SEQUELA
C2977863|T037|S32.591B|ICD10CM|OTHER SPECIFIED FRACTURE OF RIGHT PUBIS, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF RIGHT PUBIS, INIT ENCNTR FOR OPEN FRACTURE
C2857891|T037|S72.335B|ICD10CM|NONDISPLACED OBLIQUE FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP OBLIQUE FX SHAFT OF L FEMR, INIT FOR OPN FX TYPE I/2
C2977862|T037|S32.591A|ICD10CM|OTHER SPECIFIED FRACTURE OF RIGHT PUBIS, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF RIGHT PUBIS, INIT ENCNTR FOR CLOSED FRACTURE
C4270220|T046|T83.032A|ICD10CM|LEAKAGE OF NEPHROSTOMY CATHETER, INITIAL ENCOUNTER|LEAKAGE OF NEPHROSTOMY CATHETER, INITIAL ENCOUNTER
C2843271|T037|S48.011S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT RIGHT SHOULDER JOINT, SEQUELA|COMPLETE TRAUMATIC AMPUTATION AT R SHOULDER JT, SEQUELA
C2832192|T037|S06.333S|ICD10CM|CONTUSION AND LACERATION OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, SEQUELA|CONTUS/LAC CEREB, W LOC OF 1-5 HRS 59 MIN, SEQUELA
C2857892|T037|S72.335C|ICD10CM|NONDISPLACED OBLIQUE FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP OBLIQUE FX SHAFT OF L FEMR, 7THC
C2833369|T037|S12.290B|ICD10CM|OTHER DISPLACED FRACTURE OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH DISP FX OF THIRD CERVICAL VERTEBRA, INIT FOR OPN FX
C2860046|T037|S78.929S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED HIP AND THIGH, LEVEL UNSPECIFIED, SEQUELA|PARTIAL TRAUM AMP OF UNSP HIP AND THIGH, LEVEL UNSP, SEQUELA
C0348464|T046|E31.8|DMDICD10|OTHER POLYGLANDULAR DYSFUNCTION|SONSTIGE POLYGLANDULAERE DYSFUNKTION
C2878406|T037|T43.222A|ICD10CM|POISONING BY SELECTIVE SEROTONIN REUPTAKE INHIBITORS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY SLCTV SEROTONIN REUPTAKE INHIBTR, SELF-HARM, INIT
C2832190|T037|S06.333A|ICD10CM|CONTUSION AND LACERATION OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|CONTUS/LAC CEREB, W LOC OF 1-5 HRS 59 MIN, INIT
C2843269|T037|S48.011A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT RIGHT SHOULDER JOINT, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION AT RIGHT SHOULDER JOINT, INIT
C2879338|T037|T45.8X2S|ICD10CM|POISONING BY OTHER PRIMARILY SYSTEMIC AND HEMATOLOGICAL AGENTS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY OTH PRIM SYS AND HEMATOLOG AGENTS, SLF-HRM, SEQUELA
C4270431|T046|T83.82XA|ICD10CM|FIBROSIS DUE TO GENITOURINARY PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|FIBROSIS DUE TO GENITOURINARY PROSTH DEV/GRFT, INIT
C2890838|T037|T84.612A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL FIXATION DEVICE OF RIGHT RADIUS, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INT FIX OF RIGHT RADIUS, INIT
C0153658|T191|C75.9|DMDICD10|MALIGNANT NEOPLASM OF ENDOCRINE GLAND, UNSPECIFIED|BOESARTIGE NEUBILDUNG: ENDOKRINE DRUESE, NICHT NAEHER BEZEICHNET
C0348378|T191|C75.8|DMDICD10|MALIGNANT NEOPLASM WITH PLURIGLANDULAR INVOLVEMENT, UNSPECIFIED|BOESARTIGE NEUBILDUNG: BETEILIGUNG MEHRERER ENDOKRINER DRUESEN, NICHT NAEHER BEZEICHNET
C0496842|T191|C75.1|DMDICD10|MALIGNANT NEOPLASM OF PITUITARY GLAND|BOESARTIGE NEUBILDUNG: HYPOPHYSE
C0153653|T191|C75.0|DMDICD10|MALIGNANT NEOPLASM OF PARATHYROID GLAND|BOESARTIGE NEUBILDUNG: NEBENSCHILDDRUESE
C0153655|T191|C75.3|DMDICD10|MALIGNANT NEOPLASM OF PINEAL GLAND|BOESARTIGE NEUBILDUNG: EPIPHYSE [GLANDULA PINEALIS] [ZIRBELDRUESE]
C0496843|T191|C75.2|DMDICD10|MALIGNANT NEOPLASM OF CRANIOPHARYNGEAL DUCT|BOESARTIGE NEUBILDUNG: DUCTUS CRANIOPHARYNGEALIS
C2521753|T060|C755|ICD10PCS|MALIGNANT NEOPLASM OF AORTIC BODY AND OTHER PARAGANGLIA|NUCLEAR MEDICINE @ LYMPHATIC AND HEMATOLOGIC SYSTEM @ NONIMAGING NUCLEAR MEDICINE PROBE @ LYMPHATICS, HEAD AND NECK
C0153656|T191|C75.4|DMDICD10|MALIGNANT NEOPLASM OF CAROTID BODY|BOESARTIGE NEUBILDUNG: GLOMUS CAROTICUM
C2883408|T037|T49.5X2S|ICD10CM|POISONING BY OPHTHALMOLOGICAL DRUGS AND PREPARATIONS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OPTH DRUGS AND PREPARATIONS, SELF-HARM, SEQUELA
C0085860|T047||ICD10CM|AUTOIMMUNE POLYGLANDULAR FAILURE
C2883048|T047|I75.023|ICD10CM|ATHEROEMBOLISM OF BILATERAL LOWER EXTREMITIES|ATHEROEMBOLISM OF BILATERAL LOWER EXTREMITIES
C2883047|T047|I75.022|ICD10CM|ATHEROEMBOLISM OF LEFT LOWER EXTREMITY|ATHEROEMBOLISM OF LEFT LOWER EXTREMITY
C2883046|T047|I75.021|ICD10CM|ATHEROEMBOLISM OF RIGHT LOWER EXTREMITY|ATHEROEMBOLISM OF RIGHT LOWER EXTREMITY
C2883381|T037|T49.4X2A|ICD10CM|POISONING BY KERATOLYTICS, KERATOPLASTICS, AND OTHER HAIR TREATMENT DRUGS AND PREPARATIONS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY KERATOLYT/KERATPLST/HAIR TRMT DRUG, SELF-HARM, INIT
C2835183|T037|S22.009B|ICD10CM|UNSPECIFIED FRACTURE OF UNSPECIFIED THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF UNSP THORACIC VERTEBRA, INIT FOR OPN FX
C2883049|T047|I75.029|ICD10CM|ATHEROEMBOLISM OF UNSPECIFIED LOWER EXTREMITY|ATHEROEMBOLISM OF UNSPECIFIED LOWER EXTREMITY
C2883406|T037|T49.5X2A|ICD10CM|POISONING BY OPHTHALMOLOGICAL DRUGS AND PREPARATIONS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OPTH DRUGS AND PREPARATIONS, SELF-HARM, INIT
C2883383|T037|T49.4X2S|ICD10CM|POISONING BY KERATOLYTICS, KERATOPLASTICS, AND OTHER HAIR TREATMENT DRUGS AND PREPARATIONS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY KERATOLYT/KERATPLST/HAIR TRMT DRUG, SLF-HRM, SQLA
C2882671|T047|I69.952|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING LEFT DOMINANT SIDE|HEMIPLGA FOL UNSP CEREBVASC DISEASE AFF LEFT DOMINANT SIDE
C4268481|T047|I63.313|ICD10CM|CEREBRAL INFARCTION DUE TO THROMBOSIS OF BILATERAL MIDDLE CEREBRAL ARTERIES|CEREBRAL INFRC DUE TO THOMBOS OF BI MIDDLE CEREBRAL ARTERIES
C2896499|T046|M80.019A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, UNSPECIFIED SHOULDER, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FX, UNSP SHOULDER, INIT
C2888589|T047|L89.812|ICD10CM|PRESSURE ULCER OF HEAD, STAGE 2|PRESSURE ULCER OF HEAD, STAGE 2
C2888592|T047|L89.813|ICD10CM|PRESSURE ULCER OF HEAD, STAGE 3|PRESSURE ULCER OF HEAD, STAGE 3
C2888583|T047||ICD10CM|PRESSURE ULCER OF HEAD, UNSTAGEABLE
C2888586|T047|L89.811|ICD10CM|PRESSURE ULCER OF HEAD, STAGE 1|PRESSURE ULCER OF HEAD, STAGE 1
C2888595|T047|L89.814|ICD10CM|PRESSURE ULCER OF HEAD, STAGE 4|PRESSURE ULCER OF HEAD, STAGE 4
C2895176|T047|M32.9|ICD10CM|SYSTEMIC LUPUS ERYTHEMATOSUS, UNSPECIFIED|SYSTEMIC LUPUS ERYTHEMATOSUS WITHOUT ORGAN INVOLVEMENT
C2888598|T047|L89.819|ICD10CM|PRESSURE ULCER OF HEAD, UNSPECIFIED STAGE|PRESSURE ULCER OF HEAD, UNSPECIFIED STAGE
C0263591|T046|M32.0|DMDICD10|DRUG-INDUCED SYSTEMIC LUPUS ERYTHEMATOSUS|ARZNEIMITTELINDUZIERTER SYSTEMISCHER LUPUS ERYTHEMATODES
C2873807|T047|D69.42|ICD10CM|CONGENITAL AND HEREDITARY THROMBOCYTOPENIA PURPURA|CONGENITAL AND HEREDITARY THROMBOCYTOPENIA PURPURA
C0272126|T047|D69.41|ICD10CM|EVANS SYNDROME|EVANS SYNDROME
C4270235|T046|T83.091A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INDWELLING URETHRAL CATHETER, INITIAL ENCOUNTER|MECH COMPL OF INDWELLING URETHRAL CATHETER, INIT
C2833570|T037|S12.590B|ICD10CM|OTHER DISPLACED FRACTURE OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH DISP FX OF SIXTH CERVICAL VERTEBRA, INIT FOR OPN FX
C2833569|T037|S12.590A|ICD10CM|OTHER DISPLACED FRACTURE OF SIXTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH DISP FX OF SIXTH CERVICAL VERTEBRA, INIT FOR CLOS FX
C1260901|T047|D69.49|ICD10CM|OTHER PRIMARY THROMBOCYTOPENIA|MEGAKARYOCYTIC HYPOPLASIA
C2882674|T047|I69.959|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING UNSPECIFIED SIDE|HEMIPLGA FOLLOWING UNSP CEREBVASC DISEASE AFF UNSP SIDE
C2835772|T037|S24.109A|ICD10CM|UNSPECIFIED INJURY AT UNSPECIFIED LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY AT UNSP LEVEL OF THORACIC SPINAL CORD, INIT
C2891302|T046||ICD10CM|INTESTINE TRANSPLANT INFECTION
C2891301|T037|T86.851|ICD10CM|INTESTINE TRANSPLANT FAILURE|INTESTINE TRANSPLANT FAILURE
C1141940|T046||ICD10CM|INTESTINE TRANSPLANT REJECTION
C2874119|T047|E11.630|ICD10CM|TYPE 2 DIABETES MELLITUS WITH PERIODONTAL DISEASE|TYPE 2 DIABETES MELLITUS WITH PERIODONTAL DISEASE
C2891304|T037|T86.859|ICD10CM|UNSPECIFIED COMPLICATION OF INTESTINE TRANSPLANT|UNSPECIFIED COMPLICATION OF INTESTINE TRANSPLANT
C2891303|T037|T86.858|ICD10CM|OTHER COMPLICATIONS OF INTESTINE TRANSPLANT|OTHER COMPLICATIONS OF INTESTINE TRANSPLANT
C2874120|T047|E11.638|ICD10CM|TYPE 2 DIABETES MELLITUS WITH OTHER ORAL COMPLICATIONS|TYPE 2 DIABETES MELLITUS WITH OTHER ORAL COMPLICATIONS
C2883096|T047|I82.419|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED FEMORAL VEIN|ACUTE EMBOLISM AND THROMBOSIS OF UNSPECIFIED FEMORAL VEIN
C4268257|T048|F15.288|ICD10CM|OTHER STIMULANT DEPENDENCE WITH OTHER STIMULANT-INDUCED DISORDER|AMPHETAMINE OR OTHER STIMULANT USE DISORDER, SEVERE, WITH AMPHETAMINE OR OTHER STIMULANT INDUCED OBSESSIVE COMPULSIVE OR RELATED DISORDER
C4270363|T046|T83.69XA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO OTHER PROSTHETIC DEVICE, IMPLANT AND GRAFT IN GENITAL TRACT, INITIAL ENCOUNTER|I/I REACT D/T OTHER PROSTH DEV/GRFT IN GENITAL TRACT, INIT
C2874657|T048|F15.280|ICD10CM|OTHER STIMULANT DEPENDENCE WITH STIMULANT-INDUCED ANXIETY DISORDER|OTH STIMULANT DEPENDENCE W STIM-INDUCE ANXIETY DISORDER
C2874658|T048|F15.281|ICD10CM|OTHER STIMULANT DEPENDENCE WITH STIMULANT-INDUCED SEXUAL DYSFUNCTION|OTH STIMULANT DEPENDENCE W STIM-INDUCE SEXUAL DYSFUNCTION
C2874659|T048|F15.282|ICD10CM|OTHER STIMULANT DEPENDENCE WITH STIMULANT-INDUCED SLEEP DISORDER|OTH STIMULANT DEPENDENCE W STIMULANT-INDUCED SLEEP DISORDER
C2875385|T047|G95.11|ICD10CM|ACUTE INFARCTION OF SPINAL CORD (EMBOLIC) (NONEMBOLIC)|ACUTE INFARCTION OF SPINAL CORD (EMBOLIC) (NONEMBOLIC)
C2838628|T037|S34.104A|ICD10CM|UNSPECIFIED INJURY TO L4 LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|UNSP INJURY TO L4 LEVEL OF LUMBAR SPINAL CORD, INIT ENCNTR
C2838630|T037|S34.104S|ICD10CM|UNSPECIFIED INJURY TO L4 LEVEL OF LUMBAR SPINAL CORD, SEQUELA|UNSP INJURY TO L4 LEVEL OF LUMBAR SPINAL CORD, SEQUELA
C2859999|T037|S78.111S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN RIGHT HIP AND KNEE, SEQUELA|COMPLETE TRAUMATIC AMP AT LEVEL BETW R HIP AND KNEE, SEQUELA
C2883094|T047|I82.412|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF LEFT FEMORAL VEIN|ACUTE EMBOLISM AND THROMBOSIS OF LEFT FEMORAL VEIN
C4270391|T046|T83.719A|ICD10CM|EROSION OF OTHER PROSTHETIC MATERIALS TO SURROUNDING ORGAN OR TISSUE, INITIAL ENCOUNTER|EROSION OF OTHER PROSTH MATERIALS TO SURRND ORG/TISS, INIT
C2875387|T047|G95.19|ICD10CM|OTHER VASCULAR MYELOPATHIES|OTHER VASCULAR MYELOPATHIES
C2857599|T037|S72.23XB|ICD10CM|DISPLACED SUBTROCHANTERIC FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPLACED SUBTROCHNT FX UNSP FEMUR, INIT FOR OPN FX TYPE I/2
C2888539|T047|L89.603|ICD10CM|PRESSURE ULCER OF UNSPECIFIED HEEL, STAGE 3|PRESSURE ULCER OF UNSPECIFIED HEEL, STAGE 3
C2857598|T037|S72.23XA|ICD10CM|DISPLACED SUBTROCHANTERIC FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED SUBTROCHANTERIC FRACTURE OF UNSP FEMUR, INIT
C2879821|T037|T47.6X2A|ICD10CM|POISONING BY ANTIDIARRHEAL DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ANTIDIARRHEAL DRUGS, SELF-HARM, INIT
C2888533|T047|L89.601|ICD10CM|PRESSURE ULCER OF UNSPECIFIED HEEL, STAGE 1|PRESSURE ULCER OF UNSPECIFIED HEEL, STAGE 1
C2859114|T037|S72.92XB|ICD10CM|UNSPECIFIED FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP FRACTURE OF LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C2888530|T047|L89.600|ICD10CM|PRESSURE ULCER OF UNSPECIFIED HEEL, UNSTAGEABLE|PRESSURE ULCER OF UNSPECIFIED HEEL, UNSTAGEABLE
C2888254|T047|L89.100|ICD10CM|PRESSURE ULCER OF UNSPECIFIED PART OF BACK, UNSTAGEABLE|PRESSURE ULCER OF UNSPECIFIED PART OF BACK, UNSTAGEABLE
C2888257|T047|L89.101|ICD10CM|PRESSURE ULCER OF UNSPECIFIED PART OF BACK, STAGE 1|PRESSURE ULCER OF UNSPECIFIED PART OF BACK, STAGE 1
C2888260|T047|L89.102|ICD10CM|PRESSURE ULCER OF UNSPECIFIED PART OF BACK, STAGE 2|PRESSURE ULCER OF UNSPECIFIED PART OF BACK, STAGE 2
C2888263|T047|L89.103|ICD10CM|PRESSURE ULCER OF UNSPECIFIED PART OF BACK, STAGE 3|PRESSURE ULCER OF UNSPECIFIED PART OF BACK, STAGE 3
C2888266|T047|L89.104|ICD10CM|PRESSURE ULCER OF UNSPECIFIED PART OF BACK, STAGE 4|PRESSURE ULCER OF UNSPECIFIED PART OF BACK, STAGE 4
C2837978|T191|C40.32|ICD10CM|MALIGNANT NEOPLASM OF SHORT BONES OF LEFT LOWER LIMB|MALIGNANT NEOPLASM OF SHORT BONES OF LEFT LOWER LIMB
C2837977|T191|C40.31|ICD10CM|MALIGNANT NEOPLASM OF SHORT BONES OF RIGHT LOWER LIMB|MALIGNANT NEOPLASM OF SHORT BONES OF RIGHT LOWER LIMB
C2837976|T191|C40.30|ICD10CM|MALIGNANT NEOPLASM OF SHORT BONES OF UNSPECIFIED LOWER LIMB|MALIGNANT NEOPLASM OF SHORT BONES OF UNSPECIFIED LOWER LIMB
C2888269|T047|L89.109|ICD10CM|PRESSURE ULCER OF UNSPECIFIED PART OF BACK, UNSPECIFIED STAGE|PRESSURE ULCER OF UNSP PART OF BACK, UNSPECIFIED STAGE
C2900540|T046|M80.869A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, UNSPECIFIED LOWER LEG, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, UNSP LOWER LEG, INIT
C2882861|T047|I70.503|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, BILATERAL LEGS|UNSP ATHSCL NONAUT BIO BYPASS OF THE EXTRM, BILATERAL LEGS
C2882860|T047|I70.502|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, LEFT LEG|UNSP ATHSCL NONAUT BIO BYPASS OF THE EXTREMITIES, LEFT LEG
C2882859|T047|I70.501|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, RIGHT LEG|UNSP ATHSCL NONAUT BIO BYPASS OF THE EXTREMITIES, RIGHT LEG
C2882863|T047|I70.509|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, UNSPECIFIED EXTREMITY|UNSP ATHSCL NONAUT BIO BYPASS OF THE EXTRM, UNSP EXTREMITY
C2882862|T047|I70.508|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES, OTHER EXTREMITY|UNSP ATHSCL NONAUT BIO BYPASS OF THE EXTRM, OTH EXTREMITY
C0342498|T046|E27.5|ICD10CM|ADRENOMEDULLARY HYPERFUNCTION|ADRENOMEDULLARY HYPERPLASIA
C2837466|T037|S32.008A|ICD10CM|OTHER FRACTURE OF UNSPECIFIED LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF UNSP LUMBAR VERTEBRA, INIT FOR CLOS FX
C2874195|T047|E27.0|ICD10CM|OTHER ADRENOCORTICAL OVERACTIVITY|OVERPRODUCTION OF ACTH, NOT ASSOCIATED WITH CUSHING'S DISEASE
C0271737|T047|E27.1|ICD10CM|PRIMARY ADRENOCORTICAL INSUFFICIENCY|AUTOIMMUNE ADRENALITIS
C0151467|T047|E27.2|DMDICD10|ADDISONIAN CRISIS|ADDISON-KRISE
C0348943|T046|E27.3|DMDICD10|DRUG-INDUCED ADRENOCORTICAL INSUFFICIENCY|ARZNEIMITTELINDUZIERTE NEBENNIERENRINDENINSUFFIZIENZ
C0271749|T047|E27.8|ICD10CM|OTHER SPECIFIED DISORDERS OF ADRENAL GLAND|ABNORMALITY OF CORTISOL-BINDING GLOBULIN
C0001621|T047|E27.9|DMDICD10|DISORDER OF ADRENAL GLAND, UNSPECIFIED|KRANKHEIT DER NEBENNIERE, NICHT NAEHER BEZEICHNET
C2831453|T037|S02.19XA|ICD10CM|OTHER FRACTURE OF BASE OF SKULL, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF BASE OF SKULL, INIT FOR CLOS FX
C2831454|T037|S02.19XB|ICD10CM|OTHER FRACTURE OF BASE OF SKULL, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF BASE OF SKULL, INIT ENCNTR FOR OPEN FRACTURE
C2865563|T037|S88.129A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, UNSPECIFIED LOWER LEG, INITIAL ENCOUNTER|PART TRAUM AMP AT LEV BETW KNEE AND ANKL, UNSP LOW LEG, INIT
C2900889|T046|M84.421A|ICD10CM|PATHOLOGICAL FRACTURE, RIGHT HUMERUS, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, RIGHT HUMERUS, INIT FOR FX
C2865564|T037|S88.129D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, UNSPECIFIED LOWER LEG, SUBSEQUENT ENCOUNTER|PART TRAUM AMP AT LEV BETW KNEE AND ANKL, UNSP LOW LEG, SUBS
C2882747|T047|I70.302|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, LEFT LEG|UNSP ATHSCL UNSP TYPE BYPASS OF THE EXTREMITIES, LEFT LEG
C2888746|T047|L97.819|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF RIGHT LOWER LEG WITH UNSPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OTH PRT R LOW LEG W UNSP SEVERITY
C4509325|T047|L97.818|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF RIGHT LOWER LEG WITH OTHER SPECIFIED SEVERITY|NON-PRS CHRONIC ULCER OTH PRT R LOW LEG WITH OTH SEVERITY
C4509323|T047|L97.815|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF RIGHT LOWER LEG WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OTH PRT R LOW LEG W MSL INVL W/O EVD OF NECR
C2888745|T047|L97.814|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF RIGHT LOWER LEG WITH NECROSIS OF BONE|NON-PRS CHRONIC ULCER OTH PRT R LOW LEG W NECROSIS OF BONE
C4509324|T047|L97.816|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF RIGHT LOWER LEG WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OTH PRT R LOW LEG W BNE INVL W/O EVD OF NECR
C2888742|T047|L97.811|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF RIGHT LOWER LEG LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHR ULCER OTH PRT R LOW LEG LIMITED TO BRKDWN SKIN
C2888744|T047|L97.813|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF RIGHT LOWER LEG WITH NECROSIS OF MUSCLE|NON-PRS CHRONIC ULCER OTH PRT R LOW LEG W NECROSIS OF MUSCLE
C2888743|T047|L97.812|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF RIGHT LOWER LEG WITH FAT LAYER EXPOSED|NON-PRS CHRONIC ULCER OTH PRT R LOW LEG W FAT LAYER EXPOSED
C2865529|T037|S88.021A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT KNEE LEVEL, RIGHT LOWER LEG, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION AT KNEE LEVEL, R LOW LEG, INIT
C4270808|T047|H40.1121|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, LEFT EYE, MILD STAGE|PRIMARY OPEN-ANGLE GLAUCOMA, LEFT EYE, MILD STAGE
C4269270|T037|S02.112S|ICD10CM|TYPE III OCCIPITAL CONDYLE FRACTURE, UNSPECIFIED SIDE, SEQUELA|TYPE III OCCIPITAL CONDYLE FRACTURE, UNSP SIDE, SEQUELA
C2865531|T037|S88.021S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT KNEE LEVEL, RIGHT LOWER LEG, SEQUELA|PARTIAL TRAUMATIC AMP AT KNEE LEVEL, R LOW LEG, SEQUELA
C4268149|T047|E13.3511|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|OTH DIAB WITH PROLIF DIAB RTNOP WITH MACULAR EDEMA, R EYE
C4268151|T047|E13.3513|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|OTH DIAB WITH PROLIF DIABETIC RTNOP WITH MACULAR EDEMA, BI
C4268150|T047|E13.3512|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, LEFT EYE|OTH DIAB WITH PROLIF DIAB RTNOP WITH MACULAR EDEMA, LEFT EYE
C4269266|T037|S02.112B|ICD10CM|TYPE III OCCIPITAL CONDYLE FRACTURE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|TYPE III OCCIPITAL CONDYLE FRACTURE, UNSPECIFIED SIDE, 7THB
C4269265|T037|S02.112A|ICD10CM|TYPE III OCCIPITAL CONDYLE FRACTURE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE III OCCIPITAL CONDYLE FRACTURE, UNSPECIFIED SIDE, INIT
C4268152|T047|E13.3519|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH PROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|OTH DIAB WITH PROLIF DIABETIC RTNOP WITH MACULAR EDEMA, UNSP
C2832344|T037|S06.369S|ICD10CM|TRAUMATIC HEMORRHAGE OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|TRAUM HEMOR CEREB, W LOC OF UNSP DURATION, SEQUELA
C2859190|T037|S73.022A|ICD10CM|OBTURATOR SUBLUXATION OF LEFT HIP, INITIAL ENCOUNTER|OBTURATOR SUBLUXATION OF LEFT HIP, INITIAL ENCOUNTER
C4269571|T037|S02.80XS|ICD10CM|FRACTURE OF OTHER SPECIFIED SKULL AND FACIAL BONES, UNSPECIFIED SIDE, SEQUELA|FX OTH SKULL AND FACIAL BONES, UNSPECIFIED SIDE, SEQUELA
C2838509|T037|S32.89XB|ICD10CM|FRACTURE OF OTHER PARTS OF PELVIS, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF OTH PARTS OF PELVIS, INIT FOR OPN FX
C2832342|T037|S06.369A|ICD10CM|TRAUMATIC HEMORRHAGE OF CEREBRUM, UNSPECIFIED, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|TRAUM HEMOR CEREB, W LOC OF UNSP DURATION, INIT
C2873877|T047|E05.90|ICD10CM|THYROTOXICOSIS, UNSPECIFIED WITHOUT THYROTOXIC CRISIS OR STORM|THYROTOXICOSIS, UNSP WITHOUT THYROTOXIC CRISIS OR STORM
C2873878|T047|E05.91|ICD10CM|THYROTOXICOSIS, UNSPECIFIED WITH THYROTOXIC CRISIS OR STORM|THYROTOXICOSIS, UNSPECIFIED WITH THYROTOXIC CRISIS OR STORM
C2878254|T037|T42.8X2S|ICD10CM|POISONING BY ANTIPARKINSONISM DRUGS AND OTHER CENTRAL MUSCLE-TONE DEPRESSANTS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY ANTIPARKNS DRUG/CENTR MUSC-TONE DEPR, SLF-HRM, SQLA
C2833980|T037|S14.137A|ICD10CM|ANTERIOR CORD SYNDROME AT C7 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|ANTERIOR CORD SYNDROME AT C7, INIT
C2838508|T037|S32.89XA|ICD10CM|FRACTURE OF OTHER PARTS OF PELVIS, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF OTH PARTS OF PELVIS, INIT FOR CLOS FX
C2902905|T047|N05.9|ICD10CM|UNSPECIFIED NEPHRITIC SYNDROME WITH UNSPECIFIED MORPHOLOGIC CHANGES|UNSP NEPHRITIC SYNDROME WITH UNSPECIFIED MORPHOLOGIC CHANGES
C2876206|T037|T32.64|ICD10CM|CORROSIONS INVOLVING 60-69% OF BODY SURFACE WITH 40-49% THIRD DEGREE CORROSION|CORROS 60-69% OF BODY SURFACE W 40-49% THIRD DEGREE CORROS
C2889624|T047|M08.879|ICD10CM|OTHER JUVENILE ARTHRITIS, UNSPECIFIED ANKLE AND FOOT|OTHER JUVENILE ARTHRITIS, UNSPECIFIED ANKLE AND FOOT
C2876208|T037|T32.66|ICD10CM|CORROSIONS INVOLVING 60-69% OF BODY SURFACE WITH 60-69% THIRD DEGREE CORROSION|CORROS 60-69% OF BODY SURFACE W 60-69% THIRD DEGREE CORROS
C4268084|T047|E11.3411|ICD10CM|TYPE 2 DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|TYPE 2 DIAB WITH SEVERE NONP RTNOP WITH MACULAR EDEMA, R EYE
C2838022|T037|S32.413B|ICD10CM|DISPLACED FRACTURE OF ANTERIOR WALL OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISP FX OF ANTERIOR WALL OF UNSP ACETABULUM, INIT FOR OPN FX
C2874160|T047|E13.59|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH OTHER CIRCULATORY COMPLICATIONS|OTH DIABETES MELLITUS WITH OTHER CIRCULATORY COMPLICATIONS
C2876205|T037|T32.63|ICD10CM|CORROSIONS INVOLVING 60-69% OF BODY SURFACE WITH 30-39% THIRD DEGREE CORROSION|CORROS 60-69% OF BODY SURFACE W 30-39% THIRD DEGREE CORROS
C2889622|T047|M08.871|ICD10CM|OTHER JUVENILE ARTHRITIS, RIGHT ANKLE AND FOOT|OTHER JUVENILE ARTHRITIS, RIGHT ANKLE AND FOOT
C2889623|T047|M08.872|ICD10CM|OTHER JUVENILE ARTHRITIS, LEFT ANKLE AND FOOT|OTHER JUVENILE ARTHRITIS, LEFT ANKLE AND FOOT
C2886738|T037|T79.6XXA|ICD10CM|TRAUMATIC ISCHEMIA OF MUSCLE, INITIAL ENCOUNTER|TRAUMATIC ISCHEMIA OF MUSCLE, INITIAL ENCOUNTER
C2874159|T047|E13.52|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC PERIPHERAL ANGIOPATHY WITH GANGRENE|OTH DIABETES W DIABETIC PERIPHERAL ANGIOPATHY W GANGRENE
C2874157|T047|E13.51|ICD10CM|OTHER SPECIFIED DIABETES MELLITUS WITH DIABETIC PERIPHERAL ANGIOPATHY WITHOUT GANGRENE|OTH DIABETES W DIABETIC PERIPHERAL ANGIOPATHY W/O GANGRENE
C4048705|T047|E72.19|ICD10CM|OTHER DISORDERS OF SULFUR-BEARING AMINO-ACID METABOLISM|METHIONINEMIA
C0268613|T047|E72.10|ICD10CM|DISORDERS OF SULFUR-BEARING AMINO-ACID METABOLISM, UNSPECIFIED|DISORDERS OF SULFUR-BEARING AMINO-ACID METABOLISM, UNSPECIFIED
C0019880|T047|E72.11|ICD10CM|HOMOCYSTINURIA|CYSTATHIONINE SYNTHASE DEFICIENCY
C1856061|T047|E72.12|ICD10CM|METHYLENETETRAHYDROFOLATE REDUCTASE DEFICIENCY|METHYLENETETRAHYDROFOLATE REDUCTASE DEFICIENCY
C2889367|T047|M05.832|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT WRIST|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF LEFT WRIST
C2889366|T047|M05.831|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT WRIST|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF RIGHT WRIST
C2833383|T037|S12.300A|ICD10CM|UNSPECIFIED DISPLACED FRACTURE OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP DISP FX OF FOURTH CERVICAL VERTEBRA, INIT FOR CLOS FX
C2860045|T037|S78.929D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED HIP AND THIGH, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|PARTIAL TRAUM AMP OF UNSP HIP AND THIGH, LEVEL UNSP, SUBS
C2889368|T047|M05.839|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED WRIST|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF UNSP WRIST
C0026654|T047|I67.5|DMDICD10|MOYAMOYA DISEASE|MOYAMOYA-SYNDROM
C4268087|T047|E11.3419|ICD10CM|TYPE 2 DIABETES MELLITUS WITH SEVERE NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, UNSPECIFIED EYE|TYPE 2 DIAB WITH SEVERE NONP RTNOP WITH MACULAR EDEMA, UNSP
C2832655|T037|S06.896A|ICD10CM|OTHER SPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|INTCRAN INJ W LOC >24 HR W/O RET CONSC W SURV, INIT
C2883484|T037|T49.8X2S|ICD10CM|POISONING BY OTHER TOPICAL AGENTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH TOPICAL AGENTS, SELF-HARM, SEQUELA
C4237131|T048|F42.4|ICD10CM|EXCORIATION (SKIN-PICKING) DISORDER|EXCORIATION (SKIN-PICKING) DISORDER
C2876175|T037|T31.93|ICD10CM|BURNS INVOLVING 90% OR MORE OF BODY SURFACE WITH 30-39% THIRD DEGREE BURNS|BURNS OF 90%/MORE OF BODY SURFC W 30-39% THIRD DEGREE BURNS
C2876173|T037|T31.91|ICD10CM|BURNS INVOLVING 90% OR MORE OF BODY SURFACE WITH 10-19% THIRD DEGREE BURNS|BURNS OF 90%/MORE OF BODY SURFC W 10-19% THIRD DEGREE BURNS
C2876178|T037|T31.96|ICD10CM|BURNS INVOLVING 90% OR MORE OF BODY SURFACE WITH 60-69% THIRD DEGREE BURNS|BURNS OF 90%/MORE OF BODY SURFC W 60-69% THIRD DEGREE BURNS
C2876179|T037|T31.97|ICD10CM|BURNS INVOLVING 90% OR MORE OF BODY SURFACE WITH 70-79% THIRD DEGREE BURNS|BURNS OF 90%/MORE OF BODY SURFC W 70-79% THIRD DEGREE BURNS
C0349238|T048|F42.2|DMDICD10|MIXED OBSESSIONAL THOUGHTS AND ACTS|ZWANGSGEDANKEN UND -HANDLUNGEN, GEMISCHT
C3837219|T048||ICD10CM|HOARDING DISORDER
C2832657|T037|S06.896S|ICD10CM|OTHER SPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|INTCRAN INJ W LOC >24 HR W/O RET CONSC W SURV, SEQUELA
C4269566|T037|S02.80XA|ICD10CM|FRACTURE OF OTHER SPECIFIED SKULL AND FACIAL BONES, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FX OTH SKULL AND FACIAL BONES, UNSPECIFIED SIDE, INIT
C0349239|T048|F42.8|DMDICD10|OTHER OBSESSIVE-COMPULSIVE DISORDER|SONSTIGE ZWANGSSTOERUNGEN
C0028768|T048|F42.9|DMDICD10|OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED|ZWANGSSTOERUNG, NICHT NAEHER BEZEICHNET
C2874953|T048|F45.20|ICD10CM|HYPOCHONDRIACAL DISORDER, UNSPECIFIED|HYPOCHONDRIACAL DISORDER, UNSPECIFIED
C4064938|T048|F45.21|ICD10CM|HYPOCHONDRIASIS|ILLNESS ANXIETY DISORDER
C0522182|T041|F45.22|ICD10CM|BODY DYSMORPHIC DISORDER|NOSOPHOBIA
C2884764|T037|T58.12XS|ICD10CM|TOXIC EFFECT OF CARBON MONOXIDE FROM UTILITY GAS, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF CARB MONX FROM UTILITY GAS, SLF-HRM, SEQUELA
C2874954|T048|F45.29|ICD10CM|OTHER HYPOCHONDRIACAL DISORDERS|OTHER HYPOCHONDRIACAL DISORDERS
C2845872|T191|C62.00|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED UNDESCENDED TESTIS|MALIGNANT NEOPLASM OF UNSPECIFIED UNDESCENDED TESTIS
C2882322|T046|I61.6|ICD10CM|NONTRAUMATIC INTRACEREBRAL HEMORRHAGE, MULTIPLE LOCALIZED|NONTRAUMATIC INTRACEREBRAL HEMORRHAGE, MULTIPLE LOCALIZED
C2875167|T047|G43.601|ICD10CM|PERSISTENT MIGRAINE AURA WITH CEREBRAL INFARCTION, NOT INTRACTABLE, WITH STATUS MIGRAINOSUS|PERST MIGRAINE AURA W CEREBRAL INFRC, NOT NTRCT, W STAT MIGR
C1401192|T046||ICD10CM|NONTRAUMATIC INTRACEREBRAL HEMORRHAGE IN CEREBELLUM
C2882321|T046|I61.5|ICD10CM|NONTRAUMATIC INTRACEREBRAL HEMORRHAGE, INTRAVENTRICULAR|NONTRAUMATIC INTRACEREBRAL HEMORRHAGE, INTRAVENTRICULAR
C2882320|T046|I61.2|ICD10CM|NONTRAUMATIC INTRACEREBRAL HEMORRHAGE IN HEMISPHERE, UNSPECIFIED|NONTRAUMATIC INTRACEREBRAL HEMORRHAGE IN HEMISPHERE, UNSP
C1401193|T046||ICD10CM|NONTRAUMATIC INTRACEREBRAL HEMORRHAGE IN BRAIN STEM
C2882317|T046|I61.0|ICD10CM|NONTRAUMATIC INTRACEREBRAL HEMORRHAGE IN HEMISPHERE, SUBCORTICAL|DEEP INTRACEREBRAL HEMORRHAGE (NONTRAUMATIC)
C2882319|T046|I61.1|ICD10CM|NONTRAUMATIC INTRACEREBRAL HEMORRHAGE IN HEMISPHERE, CORTICAL|SUPERFICIAL INTRACEREBRAL HEMORRHAGE (NONTRAUMATIC)
C2875168|T047|G43.609|ICD10CM|PERSISTENT MIGRAINE AURA WITH CEREBRAL INFARCTION, NOT INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|PERST MIGRAINE AURA W CEREB INFRC, NOT NTRCT, W/O STAT MIGR
C2882323|T046|I61.8|ICD10CM|OTHER NONTRAUMATIC INTRACEREBRAL HEMORRHAGE|OTHER NONTRAUMATIC INTRACEREBRAL HEMORRHAGE
C3662030|T046|I61.9|ICD10CM|NONTRAUMATIC INTRACEREBRAL HEMORRHAGE, UNSPECIFIED|NONTRAUMATIC INTRACEREBRAL HEMORRHAGE, UNSPECIFIED
C2855927|T037|S68.125S|ICD10CM|PARTIAL TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF LEFT RING FINGER, SEQUELA|PARTIAL TRAUMATIC MCP AMPUTATION OF L RNG FNGR, SEQUELA
C2890797|T037|T84.498A|ICD10CM|OTHER MECHANICAL COMPLICATION OF OTHER INTERNAL ORTHOPEDIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|MECH COMPL OF INTERNAL ORTH DEVICES, IMPLNT AND GRAFTS, INIT
C2877462|T037|T39.392A|ICD10CM|POISONING BY OTHER NONSTEROIDAL ANTI-INFLAMMATORY DRUGS [NSAID], INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY OTH NONSTEROID ANTI-INFLAM DRUGS, SELF-HARM, INIT
C2882785|T047|I70.349|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF UNSPECIFIED SITE|ATHSCL UNSP TYPE BYPASS OF THE LEFT LEG W ULCER OF UNSP SITE
C2882784|T047|I70.348|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF OTHER PART OF LOWER LEG|ATHSCL UNSP TYPE BYPASS OF LEFT LEG W ULCER OTH PRT LOW LEG
C2882783|T047|I70.345|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF OTHER PART OF FOOT|ATHSCL UNSP TYPE BYPASS OF THE LEFT LEG W ULCER OTH PRT FOOT
C2882963|T047|I70.668|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, OTHER EXTREMITY|ATHSCL NONBIOL BYPASS OF THE EXTRM W GANGRENE, OTH EXTREMITY
C2858440|T037|S72.421A|ICD10CM|DISPLACED FRACTURE OF LATERAL CONDYLE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF LATERAL CONDYLE OF RIGHT FEMUR, INIT FOR CLOS FX
C2882777|T047|I70.341|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF THIGH|ATHSCL UNSP TYPE BYPASS OF THE LEFT LEG W ULCER OF THIGH
C2882779|T047|I70.343|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF ANKLE|ATHSCL UNSP TYPE BYPASS OF THE LEFT LEG W ULCER OF ANKLE
C2882778|T047|I70.342|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF CALF|ATHSCL UNSP TYPE BYPASS OF THE LEFT LEG W ULCERATION OF CALF
C4268196|T048|F01.51|ICD10CM|VASCULAR DEMENTIA WITH BEHAVIORAL DISTURBANCE|MAJOR NEUROCOGNITIVE DISORDER WITH VIOLENT BEHAVIOR
C4268192|T048|F01.50|ICD10CM|VASCULAR DEMENTIA WITHOUT BEHAVIORAL DISTURBANCE|MAJOR NEUROCOGNITIVE DISORDER WITHOUT BEHAVIORAL DISTURBANCE
C2857788|T037|S72.325B|ICD10CM|NONDISPLACED TRANSVERSE FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP TRANSVERSE FX SHAFT OF L FEMR, 7THB
C2884400|T037|T54.3X2S|ICD10CM|TOXIC EFFECT OF CORROSIVE ALKALIS AND ALKALI-LIKE SUBSTANCES, INTENTIONAL SELF-HARM, SEQUELA|TOX EFF OF CORROSV ALKALIS & ALK-LIKE SUBSTNC, SLF-HRM, SQLA
C2857721|T037|S72.321C|ICD10CM|DISPLACED TRANSVERSE FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL TRANSVERSE FX SHAFT OF R FEMR, 7THC
C2857720|T037|S72.321B|ICD10CM|DISPLACED TRANSVERSE FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL TRANSVERSE FX SHAFT OF R FEMR, 7THB
C2857719|T037|S72.321A|ICD10CM|DISPLACED TRANSVERSE FRACTURE OF SHAFT OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED TRANSVERSE FRACTURE OF SHAFT OF RIGHT FEMUR, INIT
C0206062|T047|J84.9|DMDICD10|INTERSTITIAL PULMONARY DISEASE, UNSPECIFIED|INTERSTITIELLE LUNGENKRANKHEIT, NICHT NAEHER BEZEICHNET
C2874600|T048|F14.259|ICD10CM|COCAINE DEPENDENCE WITH COCAINE-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED|COCAINE DEPENDENCE WITH COCAINE-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED
C2874598|T048|F14.250|ICD10CM|COCAINE DEPENDENCE WITH COCAINE-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|COCAINE DEPEND W COCAINE-INDUC PSYCH DISORDER W DELUSIONS
C2874599|T048|F14.251|ICD10CM|COCAINE DEPENDENCE WITH COCAINE-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|COCAINE DEPEND W COCAINE-INDUC PSYCHOTIC DISORDER W HALLUCIN
C2884398|T037|T54.3X2A|ICD10CM|TOXIC EFFECT OF CORROSIVE ALKALIS AND ALKALI-LIKE SUBSTANCES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOX EFF OF CORROSV ALKALIS & ALK-LIKE SUBSTNC, SLF-HRM, INIT
C3665339|T047|P36|DMDICD10|BACTERIAL SEPSIS OF NEWBORN, UNSPECIFIED|BAKTERIELLE SEPSIS BEIM NEUGEBORENEN
C0477920|T047|P36.8|DMDICD10|OTHER BACTERIAL SEPSIS OF NEWBORN|SONSTIGE BAKTERIELLE SEPSIS BEIM NEUGEBORENEN
C2838666|T037|S34.121A|ICD10CM|INCOMPLETE LESION OF L1 LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|INCOMPLETE LESION OF L1 LEVEL OF LUMBAR SPINAL CORD, INIT
C2885358|T037|T63.032S|ICD10CM|TOXIC EFFECT OF TAIPAN VENOM, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF TAIPAN VENOM, INTENTIONAL SELF-HARM, SEQUELA
C2838667|T037|S34.121D|ICD10CM|INCOMPLETE LESION OF L1 LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|INCOMPLETE LESION OF L1 LEVEL OF LUMBAR SPINAL CORD, SUBS
C0495408|T047|P36.0|DMDICD10|SEPSIS OF NEWBORN DUE TO STREPTOCOCCUS, GROUP B|SEPSIS BEIM NEUGEBORENEN DURCH STREPTOKOKKEN, GRUPPE B
C4509055|T048|F13.21|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC DEPENDENCE, IN REMISSION|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE DISORDER, SEVERE, IN SUSTAINED REMISSION
C0452197|T047|P36.2|DMDICD10|SEPSIS OF NEWBORN DUE TO STAPHYLOCOCCUS AUREUS|SEPSIS BEIM NEUGEBORENEN DURCH STAPHYLOCOCCUS AUREUS
C0452199|T047|P36.5|DMDICD10|SEPSIS OF NEWBORN DUE TO ANAEROBES|SEPSIS BEIM NEUGEBORENEN DURCH ANAEROBIER
C0452198|T047|P36.4|DMDICD10|SEPSIS OF NEWBORN DUE TO ESCHERICHIA COLI|SEPSIS BEIM NEUGEBORENEN DURCH ESCHERICHIA COLI
C2838668|T037|S34.121S|ICD10CM|INCOMPLETE LESION OF L1 LEVEL OF LUMBAR SPINAL CORD, SEQUELA|INCOMPLETE LESION OF L1 LEVEL OF LUMBAR SPINAL CORD, SEQUELA
C0854456|T046|I96|ICD10CM|GANGRENE, NOT ELSEWHERE CLASSIFIED|GANGRENOUS CELLULITIS
C2865590|T037|S88.929D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED LOWER LEG, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMP OF UNSP LOWER LEG, LEVEL UNSP, SUBS
C2837944|T191|C32.0|ICD10CM|MALIGNANT NEOPLASM OF GLOTTIS|MALIGNANT NEOPLASM OF LARYNGEAL COMMISSURE (ANTERIOR)(POSTERIOR)
C3647182|T191|C32.1|ICD10CM|MALIGNANT NEOPLASM OF SUPRAGLOTTIS|MALIGNANT NEOPLASM OF POSTERIOR (LARYNGEAL) SURFACE OF EPIGLOTTIS
C0153485|T191|C32.2|DMDICD10|MALIGNANT NEOPLASM OF SUBGLOTTIS|BOESARTIGE NEUBILDUNG: SUBGLOTTIS
C0153486|T191|C32.3|DMDICD10|MALIGNANT NEOPLASM OF LARYNGEAL CARTILAGE|BOESARTIGE NEUBILDUNG: LARYNXKNORPEL
C0349040|T191|C32.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF LARYNX|BOESARTIGE NEUBILDUNG: LARYNX, MEHRERE TEILBEREICHE UEBERLAPPEND
C0007107|T191|C32.9|DMDICD10|MALIGNANT NEOPLASM OF LARYNX, UNSPECIFIED|BOESARTIGE NEUBILDUNG: LARYNX, NICHT NAEHER BEZEICHNET
C0239295|T047|B37.81|ICD10AM|CANDIDAL ESOPHAGITIS|CANDIDAL OESOPHAGITIS
C2902364|T047|M89.622|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, LEFT UPPER ARM|OSTEOPATHY AFTER POLIOMYELITIS, LEFT UPPER ARM
C2902363|T047|M89.621|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, RIGHT UPPER ARM|OSTEOPATHY AFTER POLIOMYELITIS, RIGHT UPPER ARM
C2902365|T047|M89.629|ICD10CM|OSTEOPATHY AFTER POLIOMYELITIS, UNSPECIFIED UPPER ARM|OSTEOPATHY AFTER POLIOMYELITIS, UNSPECIFIED UPPER ARM
C2902450|T047|M90.572|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, LEFT ANKLE AND FOOT|OSTEONECROSIS IN DISEASES CLASSD ELSWHR, LEFT ANKLE AND FOOT
C2890622|T037|T84.121A|ICD10CM|DISPLACEMENT OF INTERNAL FIXATION DEVICE OF LEFT HUMERUS, INITIAL ENCOUNTER|DISPLACEMENT OF INT FIX OF LEFT HUMERUS, INIT
C2857686|T037|S72.302C|ICD10CM|UNSPECIFIED FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP FX SHAFT OF LEFT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2889902|T037|T82.312A|ICD10CM|BREAKDOWN (MECHANICAL) OF FEMORAL ARTERIAL GRAFT (BYPASS), INITIAL ENCOUNTER|BREAKDOWN OF FEMORAL ARTERIAL GRAFT (BYPASS), INIT
C1318500|T047||ICD10CM|NONTOXIC GOITER, UNSPECIFIED
C0348444|T047|E04.8|DMDICD10|OTHER SPECIFIED NONTOXIC GOITER|SONSTIGE NAEHER BEZEICHNETE NICHTTOXISCHE STRUMA
C2901278|T046|M84.561A|ICD10CM|PATHOLOGICAL FRACTURE IN NEOPLASTIC DISEASE, RIGHT TIBIA, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN NEOPLASTIC DISEASE, RIGHT TIBIA, INIT
C2873863|T047|E04.2|ICD10CM|NONTOXIC MULTINODULAR GOITER|MULTINODULAR (CYSTIC) GOITER NOS
C2873862|T047|E04.1|ICD10CM|NONTOXIC SINGLE THYROID NODULE|THYROID (CYSTIC) NODULE NOS
C0342114|T047|E04.0|DMDICD10|NONTOXIC DIFFUSE GOITER|NICHTTOXISCHE DIFFUSE STRUMA
C2859984|T037|S78.021A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT RIGHT HIP JOINT, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION AT RIGHT HIP JOINT, INIT ENCNTR
C2875068|T047|G35|ICD10CM|MULTIPLE SCLEROSIS|DISSEMINATED MULTIPLE SCLEROSIS
C3264375|T046|I48.92|ICD10CM|UNSPECIFIED ATRIAL FLUTTER|UNSPECIFIED ATRIAL FLUTTER
C3264374|T046|I48.91|ICD10CM|UNSPECIFIED ATRIAL FIBRILLATION|UNSPECIFIED ATRIAL FIBRILLATION
C0031315|T047|G54.6|DMDICD10|PHANTOM LIMB SYNDROME WITH PAIN|PHANTOMSCHMERZ
C0452135|T047|G54.7|DMDICD10|PHANTOM LIMB SYNDROME WITHOUT PAIN|PHANTOMGLIED OHNE SCHMERZEN
C2845968|T191||ICD10CM|SECONDARY MALIGNANT NEOPLASM OF OTHER URINARY ORGANS
C2835276|T037|S22.032A|ICD10CM|UNSTABLE BURST FRACTURE OF THIRD THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSTABLE BURST FRACTURE OF THIRD THORACIC VERTEBRA, INIT
C2835277|T037|S22.032B|ICD10CM|UNSTABLE BURST FRACTURE OF THIRD THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSTABLE BURST FX THIRD THOR VERTEBRA, INIT FOR OPN FX
C0347011|T191|C79.11|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF BLADDER|SECONDARY MALIGNANT NEOPLASM OF BLADDER
C2845967|T191|C79.10|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF UNSPECIFIED URINARY ORGANS|SECONDARY MALIGNANT NEOPLASM OF UNSPECIFIED URINARY ORGANS
C2895190|T047|M33.29|ICD10CM|POLYMYOSITIS WITH OTHER ORGAN INVOLVEMENT|POLYMYOSITIS WITH OTHER ORGAN INVOLVEMENT
C2832095|T037|S06.310A|ICD10CM|CONTUSION AND LACERATION OF RIGHT CEREBRUM WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|CONTUS/LAC RIGHT CEREBRUM W/O LOSS OF CONSCIOUSNESS, INIT
C2890945|T037|T85.09XA|ICD10CM|OTHER MECHANICAL COMPLICATION OF VENTRICULAR INTRACRANIAL (COMMUNICATING) SHUNT, INITIAL ENCOUNTER|MECH COMPL OF VENTRICULAR INTRACRANIAL SHUNT, INIT
C2895187|T047|M33.20|ICD10CM|POLYMYOSITIS, ORGAN INVOLVEMENT UNSPECIFIED|POLYMYOSITIS, ORGAN INVOLVEMENT UNSPECIFIED
C3509000|T047||ICD10CM|POLYMYOSITIS WITH RESPIRATORY INVOLVEMENT
C2895189|T047|M33.22|ICD10CM|POLYMYOSITIS WITH MYOPATHY|POLYMYOSITIS WITH MYOPATHY
C2882962|T047|I70.663|ICD10CM|ATHEROSCLEROSIS OF NONBIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, BILATERAL LEGS|ATHSCL NONBIOL BYPASS OF THE EXTRM W GANGRENE, BI LEGS
C2349307|T191|C95.12|ICD10CM|CHRONIC LEUKEMIA OF UNSPECIFIED CELL TYPE, IN RELAPSE|CHRONIC LEUKEMIA OF UNSPECIFIED CELL TYPE, IN RELAPSE
C0686589|T191||ICD10AM|CHRONIC LEUKEMIA OF UNSPECIFIED CELL TYPE, IN REMISSION
C2861646|T191|C95.10|ICD10CM|CHRONIC LEUKEMIA OF UNSPECIFIED CELL TYPE NOT HAVING ACHIEVED REMISSION|CHRONIC LEUKEMIA OF UNSP CELL TYPE NOT ACHIEVE REMISSION
C2832097|T037|S06.310S|ICD10CM|CONTUSION AND LACERATION OF RIGHT CEREBRUM WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|CONTUS/LAC RIGHT CEREBRUM W/O LOSS OF CONSCIOUSNESS, SEQUELA
C2853793|T191|C82.08|ICD10CM|FOLLICULAR LYMPHOMA GRADE I, LYMPH NODES OF MULTIPLE SITES|FOLLICULAR LYMPHOMA GRADE I, LYMPH NODES OF MULTIPLE SITES
C2853794|T191|C82.09|ICD10CM|FOLLICULAR LYMPHOMA GRADE I, EXTRANODAL AND SOLID ORGAN SITES|FOLLICULAR LYMPHOMA GRADE I, EXTRNOD AND SOLID ORGAN SITES
C2902951|T047|N17.0|ICD10CM|ACUTE KIDNEY FAILURE WITH TUBULAR NECROSIS|ACUTE KIDNEY FAILURE WITH TUBULAR NECROSIS
C2902952|T047|N17.1|ICD10CM|ACUTE KIDNEY FAILURE WITH ACUTE CORTICAL NECROSIS|ACUTE KIDNEY FAILURE WITH ACUTE CORTICAL NECROSIS
C2853789|T191|C82.04|ICD10CM|FOLLICULAR LYMPHOMA GRADE I, LYMPH NODES OF AXILLA AND UPPER LIMB|FOLLICULAR LYMPHOMA GRADE I, NODES OF AXILLA AND UPPER LIMB
C2853790|T191|C82.05|ICD10CM|FOLLICULAR LYMPHOMA GRADE I, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|FOLICLAR LYMPH GRADE I, NODES OF ING REGION AND LOWER LIMB
C2853791|T191|C82.06|ICD10CM|FOLLICULAR LYMPHOMA GRADE I, INTRAPELVIC LYMPH NODES|FOLLICULAR LYMPHOMA GRADE I, INTRAPELVIC LYMPH NODES
C2853792|T191|C82.07|ICD10CM|FOLLICULAR LYMPHOMA GRADE I, SPLEEN|FOLLICULAR LYMPHOMA GRADE I, SPLEEN
C2853785|T191|C82.00|ICD10CM|FOLLICULAR LYMPHOMA GRADE I, UNSPECIFIED SITE|FOLLICULAR LYMPHOMA GRADE I, UNSPECIFIED SITE
C2853786|T191|C82.01|ICD10CM|FOLLICULAR LYMPHOMA GRADE I, LYMPH NODES OF HEAD, FACE, AND NECK|FOLLICULAR LYMPHOMA GRADE I, NODES OF HEAD, FACE, AND NECK
C2853787|T191|C82.02|ICD10CM|FOLLICULAR LYMPHOMA GRADE I, INTRATHORACIC LYMPH NODES|FOLLICULAR LYMPHOMA GRADE I, INTRATHORACIC LYMPH NODES
C2853788|T191|C82.03|ICD10CM|FOLLICULAR LYMPHOMA GRADE I, INTRA-ABDOMINAL LYMPH NODES|FOLLICULAR LYMPHOMA GRADE I, INTRA-ABDOMINAL LYMPH NODES
C2890918|T037|T84.86XA|ICD10CM|THROMBOSIS DUE TO INTERNAL ORTHOPEDIC PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|THROMBOSIS DUE TO INTERNAL ORTHOPEDIC PROSTH DEV/GRFT, INIT
C0236763|T048|F32.4|ICD10CM|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE, IN PARTIAL REMISSION|MAJOR DEPRESSV DISORDER, SINGLE EPISODE, IN PARTIAL REMIS
C0494397|T048|F32.0|DMDICD10|MAJOR DEPRESSIVE DISORDER, SINGLE EPISODE, MILD|LEICHTE DEPRESSIVE EPISODE
C2857532|T037|S72.145C|ICD10CM|NONDISPLACED INTERTROCHANTERIC FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP INTERTROCH FX L FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2857531|T037|S72.145B|ICD10CM|NONDISPLACED INTERTROCHANTERIC FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP INTERTROCH FX LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C2857530|T037|S72.145A|ICD10CM|NONDISPLACED INTERTROCHANTERIC FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED INTERTROCHANTERIC FRACTURE OF LEFT FEMUR, INIT
C2860082|T037|S79.012A|ICD10CM|SALTER-HARRIS TYPE I PHYSEAL FRACTURE OF UPPER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SLTR-HARIS TYPE I PHYSEAL FX UPPER END OF LEFT FEMUR, INIT
C2874101|T047|E11.44|ICD10CM|TYPE 2 DIABETES MELLITUS WITH DIABETIC AMYOTROPHY|TYPE 2 DIABETES MELLITUS WITH DIABETIC AMYOTROPHY
C2838058|T037|S32.422B|ICD10CM|DISPLACED FRACTURE OF POSTERIOR WALL OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISP FX OF POSTERIOR WALL OF LEFT ACETAB, INIT FOR OPN FX
C2838057|T037|S32.422A|ICD10CM|DISPLACED FRACTURE OF POSTERIOR WALL OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF POSTERIOR WALL OF LEFT ACETABULUM, INIT
C2902451|T047|M90.579|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, UNSPECIFIED ANKLE AND FOOT|OSTEONECROSIS IN DISEASES CLASSD ELSWHR, UNSP ANKLE AND FOOT
C2891341|T046|T87.89|ICD10CM|OTHER COMPLICATIONS OF AMPUTATION STUMP|OTHER COMPLICATIONS OF AMPUTATION STUMP
C3263931|T037||ICD10CM|DEHISCENCE OF AMPUTATION STUMP
C2882541|T047|I69.242|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING LEFT DOMINANT SIDE|MONOPLG LOW LMB FOL OTH NTRM INTCRN HEMOR AFF LEFT DOM SIDE
C2882542|T047|I69.243|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING RIGHT NON-DOMINANT SIDE|MONOPLG LOW LMB FOL OTH NTRM INTCRN HEMOR AFF R NONDOM SIDE
C2882540|T047|I69.241|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING RIGHT DOMINANT SIDE|MONOPLG LOW LMB FOL OTH NTRM INTCRN HEMOR AFF RIGHT DOM SIDE
C2882543|T047|I69.244|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING LEFT NON-DOMINANT SIDE|MONOPLG LOW LMB FOL OTH NTRM INTCRN HEMOR AFF L NONDOM SIDE
C2882544|T047|I69.249|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING UNSPECIFIED SIDE|MONOPLG LOW LMB FOL OTH NTRM INTCRN HEMOR AFF UNSP SIDE
C2882254|T047|I42.9|ICD10CM|CARDIOMYOPATHY, UNSPECIFIED|CARDIOMYOPATHY (PRIMARY) (SECONDARY) NOS
C0348617|T047|I42.8|DMDICD10|OTHER CARDIOMYOPATHIES|SONSTIGE KARDIOMYOPATHIEN
C0700053|T019||ICD10CM|OBSTRUCTIVE HYPERTROPHIC CARDIOMYOPATHY
C0007193|T047|I42.0|DMDICD10|DILATED CARDIOMYOPATHY|DILATATIVE KARDIOMYOPATHIE
C2882252|T047||ICD10CM|ENDOMYOCARDIAL (EOSINOPHILIC) DISEASE
C0348615|T047|I42.2|DMDICD10|OTHER HYPERTROPHIC CARDIOMYOPATHY|SONSTIGE HYPERTROPHISCHE KARDIOMYOPATHIE
C0348616|T047|I42.5|DMDICD10|OTHER RESTRICTIVE CARDIOMYOPATHY|SONSTIGE RESTRIKTIVE KARDIOMYOPATHIE
C1391997|T047|I42.4|ICD10CM|ENDOCARDIAL FIBROELASTOSIS|CONGENITAL CARDIOMYOPATHY
C2882253|T047|I42.7|ICD10CM|CARDIOMYOPATHY DUE TO DRUG AND EXTERNAL AGENT|CARDIOMYOPATHY DUE TO DRUG AND EXTERNAL AGENT
C0007192|T047|I42.6|DMDICD10|ALCOHOLIC CARDIOMYOPATHY|ALKOHOLISCHE KARDIOMYOPATHIE
C2889525|T047|M08.00|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE|UNSP JUVENILE RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE
C2877150|T037|T38.6X2S|ICD10CM|POISONING BY ANTIGONADOTROPHINS, ANTIESTROGENS, ANTIANDROGENS, NOT ELSEWHERE CLASSIFIED, INTENTIONAL SELF-HARM, SEQUELA|POISN BY ANTIGONADTR/ANTIESTR/ANTIANDRG, NEC, SLF-HRM, SQLA
C2889549|T047|M08.08|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, VERTEBRAE|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, VERTEBRAE
C2889550|T047|M08.09|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, MULTIPLE SITES|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, MULTIPLE SITES
C2890699|T037|T84.213A|ICD10CM|BREAKDOWN (MECHANICAL) OF INTERNAL FIXATION DEVICE OF BONES OF FOOT AND TOES, INITIAL ENCOUNTER|BREAKDOWN OF INT FIX OF BONES OF FOOT AND TOES, INIT
C2835349|T037|S22.052B|ICD10CM|UNSTABLE BURST FRACTURE OF T5-T6 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSTABLE BURST FRACTURE OF T5-T6 VERTEBRA, INIT FOR OPN FX
C2835348|T037|S22.052A|ICD10CM|UNSTABLE BURST FRACTURE OF T5-T6 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSTABLE BURST FRACTURE OF T5-T6 VERTEBRA, INIT FOR CLOS FX
C2835828|T037|S24.143S|ICD10CM|BROWN-SEQUARD SYNDROME AT T7-T10 LEVEL OF THORACIC SPINAL CORD, SEQUELA|BROWN-SEQUARD SYNDROME AT T7-T10, SEQUELA
C2877148|T037|T38.6X2A|ICD10CM|POISONING BY ANTIGONADOTROPHINS, ANTIESTROGENS, ANTIANDROGENS, NOT ELSEWHERE CLASSIFIED, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY ANTIGONADTR/ANTIESTR/ANTIANDRG, NEC, SLF-HRM, INIT
C2835827|T037|S24.143D|ICD10CM|BROWN-SEQUARD SYNDROME AT T7-T10 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|BROWN-SEQUARD SYNDROME AT T7-T10, SUBS
C2835809|T037|S24.134A|ICD10CM|ANTERIOR CORD SYNDROME AT T11-T12 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|ANTERIOR CORD SYNDROME AT T11-T12, INIT
C2835826|T037|S24.143A|ICD10CM|BROWN-SEQUARD SYNDROME AT T7-T10 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|BROWN-SEQUARD SYNDROME AT T7-T10, INIT
C2835810|T037|S24.134D|ICD10CM|ANTERIOR CORD SYNDROME AT T11-T12 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|ANTERIOR CORD SYNDROME AT T11-T12, SUBS
C2874225|T047|E66.01|ICD10CM|MORBID (SEVERE) OBESITY DUE TO EXCESS CALORIES|MORBID (SEVERE) OBESITY DUE TO EXCESS CALORIES
C2889594|T047|M08.469|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED KNEE|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, UNSP KNEE
C2889593|T047|M08.462|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, LEFT KNEE|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, LEFT KNEE
C2889592|T047|M08.461|ICD10CM|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, RIGHT KNEE|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, RIGHT KNEE
C0494666|T047|J67|DMDICD10|HYPERSENSITIVITY PNEUMONITIS DUE TO UNSPECIFIED ORGANIC DUST|ALLERGISCHE ALVEOLITIS DURCH ORGANISCHEN STAUB
C0348697|T047|J67.8|DMDICD10|HYPERSENSITIVITY PNEUMONITIS DUE TO OTHER ORGANIC DUSTS|ALLERGISCHE ALVEOLITIS DURCH ORGANISCHE STAEUBE
C2905816|T037|X83.2XXS|ICD10CM|INTENTIONAL SELF-HARM BY EXPOSURE TO EXTREMES OF COLD, SEQUELA|SELF-HARM BY EXPOSURE TO EXTREMES OF COLD, SEQUELA
C2887474|T047|J67.1|ICD10CM|BAGASSOSIS|BAGASSE PNEUMONITIS
C2887473|T047|J67.0|ICD10CM|FARMER'S LUNG|HAYMAKER'S LUNG
C0152108|T047|J67.3|DMDICD10|SUBEROSIS|SUBEROSE
C0085931|T047||ICD10CM|BIRD FANCIER'S LUNG
C0155889|T047|J67.5|DMDICD10|MUSHROOM-WORKER'S LUNG|PILZARBEITER-LUNGE
C0155888|T047|J67.4|DMDICD10|MALTWORKER'S LUNG|MALZARBEITER-LUNGE
C2887475|T047|J67.7|ICD10CM|AIR CONDITIONER AND HUMIDIFIER LUNG|ALLERGIC ALVEOLITIS DUE TO FUNGAL, THERMOPHILIC ACTINOMYCETES AND OTHER ORGANISMS GROWING IN VENTILATION [AIR CONDITIONING] SYSTEMS
C0155890|T047|J67.6|DMDICD10|MAPLE-BARK-STRIPPER'S LUNG|AHORNRINDENSCHAELER-LUNGE
C2882637|T047|I69.864|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING LEFT NON-DOMINANT SIDE|OTH PARLYT SYND FOL OTH CEREBVASC DIS AFF LEFT NONDOM SIDE
C0393570|T047|G31.85|ICD10CM|CORTICOBASAL DEGENERATION|CORTICOBASAL DEGENERATION
C0023264|T047||ICD10CM|LEIGH'S DISEASE
C2882636|T047|I69.863|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING RIGHT NON-DOMINANT SIDE|OTH PARLYT SYND FOL OTH CEREBVASC DIS AFF RIGHT NONDOM SIDE
C0205710|T047||ICD10CM|ALPERS DISEASE
C2882639|T047|I69.869|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING UNSPECIFIED SIDE|OTH PARLYT SYNDROME FOL OTH CEREBVASC DISEASE AFF UNSP SIDE
C2842127|T191|C50.811|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF RIGHT FEMALE BREAST|MALIGNANT NEOPLASM OF OVRLP SITES OF RIGHT FEMALE BREAST
C2842128|T191|C50.812|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF LEFT FEMALE BREAST|MALIGNANT NEOPLASM OF OVRLP SITES OF LEFT FEMALE BREAST
C2833241|T037|S12.112A|ICD10CM|NONDISPLACED TYPE II DENS FRACTURE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED TYPE II DENS FRACTURE, INIT FOR CLOS FX
C3264033|T047|G43.831|ICD10CM|MENSTRUAL MIGRAINE, INTRACTABLE, WITH STATUS MIGRAINOSUS|MENSTRUAL MIGRAINE, INTRACTABLE, WITH STATUS MIGRAINOSUS
C2833242|T037|S12.112B|ICD10CM|NONDISPLACED TYPE II DENS FRACTURE, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISPLACED TYPE II DENS FRACTURE, INIT FOR OPN FX
C2842129|T191|C50.819|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF UNSPECIFIED FEMALE BREAST|MALIGNANT NEOPLASM OF OVRLP SITES OF UNSP FEMALE BREAST
C2832517|T037|S06.6X2A|ICD10CM|TRAUMATIC SUBARACHNOID HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|TRAUM SUBRAC HEM W LOSS OF CONSCIOUSNESS OF 31-59 MIN, INIT
C2890048|T037|T82.524A|ICD10CM|DISPLACEMENT OF INFUSION CATHETER, INITIAL ENCOUNTER|DISPLACEMENT OF INFUSION CATHETER, INITIAL ENCOUNTER
C3264034|T047|G43.839|ICD10CM|MENSTRUAL MIGRAINE, INTRACTABLE, WITHOUT STATUS MIGRAINOSUS|MENSTRUAL MIGRAINE, INTRACTABLE, WITHOUT STATUS MIGRAINOSUS
C2877565|T037|T40.0X2S|ICD10CM|POISONING BY OPIUM, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OPIUM, INTENTIONAL SELF-HARM, SEQUELA
C2878895|T037|T44.6X2A|ICD10CM|POISONING BY ALPHA-ADRENORECEPTOR ANTAGONISTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY ALPHA-ADRENOCPT ANTAGONISTS, SELF-HARM, INIT
C2877563|T037|T40.0X2A|ICD10CM|POISONING BY OPIUM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OPIUM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER
C2977160|T037|T87.0X9|ICD10CM|COMPLICATIONS OF REATTACHED (PART OF) UNSPECIFIED UPPER EXTREMITY|COMPLICATIONS OF REATTACHED (PART OF) UNSP UPPER EXTREMITY
C2890584|T037|T84.111A|ICD10CM|BREAKDOWN (MECHANICAL) OF INTERNAL FIXATION DEVICE OF LEFT HUMERUS, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF INT FIX OF LEFT HUMERUS, INIT
C2878897|T037|T44.6X2S|ICD10CM|POISONING BY ALPHA-ADRENORECEPTOR ANTAGONISTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY ALPHA-ADRENOCPT ANTAGONISTS, SELF-HARM, SEQUELA
C3264196|T047|H40.1220|ICD10CM|LOW-TENSION GLAUCOMA, LEFT EYE, STAGE UNSPECIFIED|LOW-TENSION GLAUCOMA, LEFT EYE, STAGE UNSPECIFIED
C2883110|T047|I82.443|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF TIBIAL VEIN, BILATERAL|ACUTE EMBOLISM AND THROMBOSIS OF TIBIAL VEIN, BILATERAL
C2883109|T047|I82.442|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF LEFT TIBIAL VEIN|ACUTE EMBOLISM AND THROMBOSIS OF LEFT TIBIAL VEIN
C2883108|T047|I82.441|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF RIGHT TIBIAL VEIN|ACUTE EMBOLISM AND THROMBOSIS OF RIGHT TIBIAL VEIN
C2859248|T037|S73.044A|ICD10CM|CENTRAL DISLOCATION OF RIGHT HIP, INITIAL ENCOUNTER|CENTRAL DISLOCATION OF RIGHT HIP, INITIAL ENCOUNTER
C2889989|T037|T82.43XS|ICD10CM|LEAKAGE OF VASCULAR DIALYSIS CATHETER, SEQUELA|LEAKAGE OF VASCULAR DIALYSIS CATHETER, SEQUELA
C2874824|T048|F19.251|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH PSYCHOACTIVE SUBSTANCE-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS|OTH PSYCHOACTV SUBSTANCE DEPEND W PSYCH DISORDER W HALLUCIN
C2874823|T048|F19.250|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH PSYCHOACTIVE SUBSTANCE-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS|OTH PSYCHOACTV SUBSTANCE DEPEND W PSYCH DISORDER W DELUSIONS
C0014518|T047|L51.2|DMDICD10|TOXIC EPIDERMAL NECROLYSIS [LYELL]|TOXISCHE EPIDERMALE NEKROLYSE [LYELL-SYNDROM]
C2349616|T047|L51.3|ICD10CM|STEVENS-JOHNSON SYNDROME-TOXIC EPIDERMAL NECROLYSIS OVERLAP SYNDROME|STEVENS-JOHNSON SYND-TOX EPDRML NECROLYSIS OVERLAP SYNDROME
C0038325|T047|L51.1|DMDICD10|STEVENS-JOHNSON SYNDROME|BULLOESES ERYTHEMA EXSUDATIVUM MULTIFORME
C2855869|T037|S68.111S|ICD10CM|COMPLETE TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF LEFT INDEX FINGER, SEQUELA|COMPLETE TRAUMATIC MCP AMPUTATION OF L IDX FNGR, SEQUELA
C2889246|T047|M05.44|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF HAND
C2855970|T037|S68.429S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED HAND AT WRIST LEVEL, SEQUELA|PARTIAL TRAUMATIC AMP OF UNSP HAND AT WRIST LEVEL, SEQUELA
C2889988|T037|T82.43XD|ICD10CM|LEAKAGE OF VASCULAR DIALYSIS CATHETER, SUBSEQUENT ENCOUNTER|LEAKAGE OF VASCULAR DIALYSIS CATHETER, SUBSEQUENT ENCOUNTER
C2889248|T047|M05.442|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT HAND|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT HAND
C2889247|T047|M05.441|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT HAND|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT HAND
C0155582|T047||ICD10CM|RHEUMATIC HEART FAILURE
C2833944|T037|S14.127D|ICD10CM|CENTRAL CORD SYNDROME AT C7 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|CENTRAL CORD SYNDROME AT C7, SUBS
C2833943|T037|S14.127A|ICD10CM|CENTRAL CORD SYNDROME AT C7 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|CENTRAL CORD SYNDROME AT C7, INIT
C2883164|T047|I82.623|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF DEEP VEINS OF UPPER EXTREMITY, BILATERAL|ACUTE EMBOLISM AND THOMBOS OF DEEP VEINS OF UP EXTREM, BI
C2883163|T047|I82.622|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF DEEP VEINS OF LEFT UPPER EXTREMITY|ACUTE EMBOLISM AND THROMBOSIS OF DEEP VEINS OF L UP EXTREM
C2883162|T047|I82.621|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF DEEP VEINS OF RIGHT UPPER EXTREMITY|ACUTE EMBOLISM AND THROMBOSIS OF DEEP VEINS OF R UP EXTREM
C2848430|T037|S58.121S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN ELBOW AND WRIST, RIGHT ARM, SEQUELA|PART TRAUM AMP AT LEV BETW ELBOW AND WRIST, RIGHT ARM, SQLA
C2856793|T037|S72.041A|ICD10CM|DISPLACED FRACTURE OF BASE OF NECK OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF BASE OF NECK OF RIGHT FEMUR, INIT FOR CLOS FX
C2883165|T047|I82.629|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF DEEP VEINS OF UNSPECIFIED UPPER EXTREMITY|ACUTE EMBOLISM AND THROMBOSIS OF DEEP VN UNSP UP EXTREM
C2856795|T037|S72.041C|ICD10CM|DISPLACED FRACTURE OF BASE OF NECK OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF BASE OF NK OF R FEMR, INIT FOR OPN FX TYPE 3A/B/C
C2843340|T037|S48.922S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT SHOULDER AND UPPER ARM, LEVEL UNSPECIFIED, SEQUELA|PARTIAL TRAUM AMP OF LEFT SHLDR/UP ARM, LEVEL UNSP, SEQUELA
C2884480|T037|T56.1X2A|ICD10CM|TOXIC EFFECT OF MERCURY AND ITS COMPOUNDS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF MERCURY AND ITS COMPOUNDS, SELF-HARM, INIT
C2889320|T047|M05.669|ICD10CM|RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF UNSP KNEE W INVOLV OF ORGANS AND SYSTEMS
C2874392|T048|F10.239|ICD10CM|ALCOHOL DEPENDENCE WITH WITHDRAWAL, UNSPECIFIED|ALCOHOL DEPENDENCE WITH WITHDRAWAL, UNSPECIFIED
C2889319|T047|M05.662|ICD10CM|RHEUMATOID ARTHRITIS OF LEFT KNEE WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF LEFT KNEE W INVOLV OF ORGANS AND SYSTEMS
C2889318|T047|M05.661|ICD10CM|RHEUMATOID ARTHRITIS OF RIGHT KNEE WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF RIGHT KNEE W INVOLV OF ORGANS AND SYSTEMS
C2874391|T048|F10.232|ICD10CM|ALCOHOL DEPENDENCE WITH WITHDRAWAL WITH PERCEPTUAL DISTURBANCE|ALCOHOL DEPENDENCE W WITHDRAWAL WITH PERCEPTUAL DISTURBANCE
C2874389|T048||ICD10CM|ALCOHOL DEPENDENCE WITH WITHDRAWAL, UNCOMPLICATED
C2874390|T048|F10.231|ICD10CM|ALCOHOL DEPENDENCE WITH WITHDRAWAL DELIRIUM|ALCOHOL DEPENDENCE WITH WITHDRAWAL DELIRIUM
C2876972|T037|T37.92XS|ICD10CM|POISONING BY UNSPECIFIED SYSTEMIC ANTI-INFECTIVE AND ANTIPARASITICS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY UNSP SYS ANTI-INFECT AND ANTIPARASTC, SLF-HRM, SQLA
C2874432|T048|F11.188|ICD10CM|OPIOID ABUSE WITH OTHER OPIOID-INDUCED DISORDER|OPIOID ABUSE WITH OTHER OPIOID-INDUCED DISORDER
C2842068|T191|C4A.61|ICD10CM|MERKEL CELL CARCINOMA OF RIGHT UPPER LIMB, INCLUDING SHOULDER|MERKEL CELL CARCINOMA OF RIGHT UPPER LIMB, INC SHOULDER
C2977925|T191|C4A.60|ICD10CM|MERKEL CELL CARCINOMA OF UNSPECIFIED UPPER LIMB, INCLUDING SHOULDER|MERKEL CELL CARCINOMA OF UNSP UPPER LIMB, INCLUDING SHOULDER
C2842069|T191|C4A.62|ICD10CM|MERKEL CELL CARCINOMA OF LEFT UPPER LIMB, INCLUDING SHOULDER|MERKEL CELL CARCINOMA OF LEFT UPPER LIMB, INCLUDING SHOULDER
C2874434|T048|F11.182|ICD10CM|OPIOID ABUSE WITH OPIOID-INDUCED SLEEP DISORDER|OPIOID ABUSE WITH OPIOID-INDUCED SLEEP DISORDER
C2874433|T048|F11.181|ICD10CM|OPIOID ABUSE WITH OPIOID-INDUCED SEXUAL DYSFUNCTION|OPIOID ABUSE WITH OPIOID-INDUCED SEXUAL DYSFUNCTION
C2876970|T037|T37.92XA|ICD10CM|POISONING BY UNSPECIFIED SYSTEMIC ANTI-INFECTIVE AND ANTIPARASITICS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY UNSP SYS ANTI-INFECT AND ANTIPARASTC, SLF-HRM, INIT
C2873773|T047|D57.81|ICD10CM|OTHER SICKLE-CELL DISORDERS WITH CRISIS, UNSPECIFIED|OTHER SICKLE-CELL DISORDERS WITH CRISIS
C2857582|T037|S72.22XB|ICD10CM|DISPLACED SUBTROCHANTERIC FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPLACED SUBTROCHNT FX LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C2857581|T037|S72.22XA|ICD10CM|DISPLACED SUBTROCHANTERIC FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED SUBTROCHANTERIC FRACTURE OF LEFT FEMUR, INIT
C0030481|T047|G04.1|DMDICD10|TROPICAL SPASTIC PARAPLEGIA|TROPISCHE SPASTISCHE PARAPLEGIE
C2873771|T047|D57.811|ICD10CM|OTHER SICKLE-CELL DISORDERS WITH ACUTE CHEST SYNDROME|OTHER SICKLE-CELL DISORDERS WITH ACUTE CHEST SYNDROME
C2873772|T047|D57.812|ICD10CM|OTHER SICKLE-CELL DISORDERS WITH SPLENIC SEQUESTRATION|OTHER SICKLE-CELL DISORDERS WITH SPLENIC SEQUESTRATION
C2882585|T047|I69.349|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING CEREBRAL INFARCTION AFFECTING UNSPECIFIED SIDE|MONOPLG LOW LMB FOLLOWING CEREBRAL INFRC AFFECTING UNSP SIDE
C2837561|T037|S32.031B|ICD10CM|STABLE BURST FRACTURE OF THIRD LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|STABLE BURST FRACTURE OF THIRD LUM VERTEBRA, INIT FOR OPN FX
C2837560|T037|S32.031A|ICD10CM|STABLE BURST FRACTURE OF THIRD LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|STABLE BURST FRACTURE OF THIRD LUMBAR VERTEBRA, INIT
C2843312|T037|S48.122A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN LEFT SHOULDER AND ELBOW, INITIAL ENCOUNTER|PARTIAL TRAUM AMP AT LEVEL BETW L SHOULDER AND ELBOW, INIT
C2848428|T037|S58.121A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN ELBOW AND WRIST, RIGHT ARM, INITIAL ENCOUNTER|PART TRAUM AMP AT LEV BETW ELBOW AND WRIST, RIGHT ARM, INIT
C2835463|T037|S22.088A|ICD10CM|OTHER FRACTURE OF T11-T12 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF T11-T12 VERTEBRA, INIT FOR CLOS FX
C2835464|T037|S22.088B|ICD10CM|OTHER FRACTURE OF T11-T12 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF T11-T12 VERTEBRA, INIT FOR OPN FX
C2879923|T037|T48.0X2S|ICD10CM|POISONING BY OXYTOCIC DRUGS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OXYTOCIC DRUGS, INTENTIONAL SELF-HARM, SEQUELA
C2890345|T037|T83.428A|ICD10CM|DISPLACEMENT OF OTHER PROSTHETIC DEVICES, IMPLANTS AND GRAFTS OF GENITAL TRACT, INITIAL ENCOUNTER|DISPLACEMENT OF PROSTH DEV/IMPLNT/GRFT OF GENITL TRCT, INIT
C4268831|T046|M97.02XA|ICD10CM|PERIPROSTHETIC FRACTURE AROUND INTERNAL PROSTHETIC LEFT HIP JOINT, INITIAL ENCOUNTER|PERIPROSTH FRACTURE AROUND INTERNAL PROSTH L HIP JT, INIT
C2858696|T037|S72.444B|ICD10CM|NONDISPLACED FRACTURE OF LOWER EPIPHYSIS (SEPARATION) OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF LOW EPIPHY (SEPARATION) OF R FEMR, 7THB
C2879921|T037|T48.0X2A|ICD10CM|POISONING BY OXYTOCIC DRUGS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OXYTOCIC DRUGS, INTENTIONAL SELF-HARM, INIT
C2875008|T048|F98.4|ICD10CM|STEREOTYPED MOVEMENT DISORDERS|STEREOTYPE/HABIT DISORDER
C2858459|T037|S72.422C|ICD10CM|DISPLACED FRACTURE OF LATERAL CONDYLE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF LATERAL CONDYLE OF L FEMR, 7THC
C4268474|T046|I16.9|ICD10CM|HYPERTENSIVE CRISIS, UNSPECIFIED|HYPERTENSIVE CRISIS, UNSPECIFIED
C2858457|T037|S72.422A|ICD10CM|DISPLACED FRACTURE OF LATERAL CONDYLE OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF LATERAL CONDYLE OF LEFT FEMUR, INIT FOR CLOS FX
C2858817|T037|S72.455B|ICD10CM|NONDISPLACED SUPRACONDYLAR FRACTURE WITHOUT INTRACONDYLAR EXTENSION OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP SUPRCNDL FX W/O INTRCNDL EXTN LOW END L FEMR, 7THB
C2845923|T191|C69.81|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF RIGHT EYE AND ADNEXA|MALIGNANT NEOPLASM OF OVRLP SITES OF RIGHT EYE AND ADNEXA
C2845922|T191|C69.80|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF UNSPECIFIED EYE AND ADNEXA|MALIGNANT NEOPLASM OF OVRLP SITES OF UNSP EYE AND ADNEXA
C2845924|T191|C69.82|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF LEFT EYE AND ADNEXA|MALIGNANT NEOPLASM OF OVRLP SITES OF LEFT EYE AND ADNEXA
C0745138|T047|I16.0|ICD10CM|HYPERTENSIVE URGENCY|HYPERTENSIVE URGENCY
C0745136|T047|I16.1|ICD10CM|HYPERTENSIVE EMERGENCY|HYPERTENSIVE EMERGENCY
C2882584|T047|I69.344|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING CEREBRAL INFARCTION AFFECTING LEFT NON-DOMINANT SIDE|MONOPLG LOW LMB FOL CEREBRAL INFRC AFF LEFT NONDOM SIDE
C2832352|T037|S06.371S|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF CEREBELLUM WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, SEQUELA|CONTUS/LAC/HEM CRBLM W LOC OF 30 MINUTES OR LESS, SEQUELA
C2869906|T037|S98.922S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT FOOT, LEVEL UNSPECIFIED, SEQUELA|PARTIAL TRAUMATIC AMP OF LEFT FOOT, LEVEL UNSP, SEQUELA
C2869905|T037|S98.922D|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT FOOT, LEVEL UNSPECIFIED, SUBSEQUENT ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF LEFT FOOT, LEVEL UNSP, SUBS
C2869904|T037|S98.922A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF LEFT FOOT, LEVEL UNSPECIFIED, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMPUTATION OF LEFT FOOT, LEVEL UNSP, INIT
C2832350|T037|S06.371A|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF CEREBELLUM WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS, INITIAL ENCOUNTER|CONTUS/LAC/HEM CRBLM W LOC OF 30 MINUTES OR LESS, INIT
C2889461|T046|M06.369|ICD10CM|RHEUMATOID NODULE, UNSPECIFIED KNEE|RHEUMATOID NODULE, UNSPECIFIED KNEE
C2889460|T046|M06.362|ICD10CM|RHEUMATOID NODULE, LEFT KNEE|RHEUMATOID NODULE, LEFT KNEE
C2889459|T046|M06.361|ICD10CM|RHEUMATOID NODULE, RIGHT KNEE|RHEUMATOID NODULE, RIGHT KNEE
C2857632|T037|S72.25XA|ICD10CM|NONDISPLACED SUBTROCHANTERIC FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED SUBTROCHANTERIC FRACTURE OF LEFT FEMUR, INIT
C4237251|T048|F11.982|ICD10CM|OPIOID USE, UNSPECIFIED WITH OPIOID-INDUCED SLEEP DISORDER|OPIOID INDUCED SLEEP DISORDER, WITHOUT USE DISORDER
C4237248|T048|F11.981|ICD10CM|OPIOID USE, UNSPECIFIED WITH OPIOID-INDUCED SEXUAL DYSFUNCTION|OPIOID INDUCED SEXUAL DYSFUNCTION, WITHOUT USE DISORDER
C2890825|T037|T84.60XA|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL FIXATION DEVICE OF UNSPECIFIED SITE, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INT FIX OF UNSP SITE, INIT
C4237242|T048|F11.988|ICD10CM|OPIOID USE, UNSPECIFIED WITH OTHER OPIOID-INDUCED DISORDER|OPIOID INDUCED ANXIETY DISORDER, WITHOUT USE DISORDER
C2857633|T037|S72.25XB|ICD10CM|NONDISPLACED SUBTROCHANTERIC FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP SUBTROCHNT FX LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C2882903|T047|I70.561|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, RIGHT LEG|ATHSCL NONAUT BIO BYPASS OF THE EXTRM W GANGRENE, RIGHT LEG
C2882905|T047|I70.563|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, BILATERAL LEGS|ATHSCL NONAUT BIO BYPASS OF THE EXTRM W GANGRENE, BI LEGS
C2882904|T047|I70.562|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, LEFT LEG|ATHSCL NONAUT BIO BYPASS OF THE EXTRM W GANGRENE, LEFT LEG
C2861674|T191|D03.51|ICD10CM|MELANOMA IN SITU OF ANAL SKIN|MELANOMA IN SITU OF ANAL SKIN
C2857684|T037|S72.302A|ICD10CM|UNSPECIFIED FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF SHAFT OF LEFT FEMUR, INIT FOR CLOS FX
C2857685|T037|S72.302B|ICD10CM|UNSPECIFIED FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|UNSP FX SHAFT OF LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C2861675|T191|D03.52|ICD10CM|MELANOMA IN SITU OF BREAST (SKIN) (SOFT TISSUE)|MELANOMA IN SITU OF BREAST (SKIN) (SOFT TISSUE)
C2882907|T047|I70.569|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, UNSPECIFIED EXTREMITY|ATHSCL NONAUT BIO BYPASS OF THE EXTRM W GANGRENE, UNSP EXTRM
C2882906|T047|I70.568|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, OTHER EXTREMITY|ATHSCL NONAUT BIO BYPASS OF THE EXTRM W GANGRENE, OTH EXTRM
C2838322|T037|S32.483A|ICD10CM|DISPLACED DOME FRACTURE OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED DOME FRACTURE OF UNSP ACETABULUM, INIT FOR CLOS FX
C2861676|T191|D03.59|ICD10CM|MELANOMA IN SITU OF OTHER PART OF TRUNK|MELANOMA IN SITU OF OTHER PART OF TRUNK
C2885075|T037|T60.4X2A|ICD10CM|TOXIC EFFECT OF RODENTICIDES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF RODENTICIDES, INTENTIONAL SELF-HARM, INIT
C2877202|T037|T38.802S|ICD10CM|POISONING BY UNSPECIFIED HORMONES AND SYNTHETIC SUBSTITUTES, INTENTIONAL SELF-HARM, SEQUELA|POISN BY UNSP HORMONES AND SYNTHETIC SUB, SELF-HARM, SEQUELA
C4269417|T037|S02.40FS|ICD10CM|ZYGOMATIC FRACTURE, LEFT SIDE, SEQUELA|ZYGOMATIC FRACTURE, LEFT SIDE, SEQUELA
C0852654|T047||ICD10CM|CONGENITAL ADRENOGENITAL DISORDERS ASSOCIATED WITH ENZYME DEFICIENCY
C0348483|T047|E70.8|DMDICD10|OTHER DISORDERS OF AROMATIC AMINO-ACID METABOLISM|SONSTIGE STOERUNGEN DES STOFFWECHSELS AROMATISCHER AMINOSAEUREN
C0342674|T047|E70|DMDICD10|DISORDER OF AROMATIC AMINO-ACID METABOLISM, UNSPECIFIED|STOERUNGEN DES STOFFWECHSELS AROMATISCHER AMINOSAEUREN
C4269413|T037|S02.40FB|ICD10CM|ZYGOMATIC FRACTURE, LEFT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|ZYGOMATIC FRACTURE, LEFT SIDE, 7THB
C0041254|T046||ICD10CM|DISORDERS OF TRYPTOPHAN METABOLISM
C1384854|T047||ICD10CM|OTHER ADRENOGENITAL DISORDERS
C0701163|T047|E25|DMDICD10|ADRENOGENITAL DISORDER, UNSPECIFIED|ADRENOGENITALE STOERUNGEN
C0751434|T047|E70.0|DMDICD10|CLASSICAL PHENYLKETONURIA|KLASSISCHE PHENYLKETONURIE
C0348482|T047|E70.1|DMDICD10|OTHER HYPERPHENYLALANINEMIAS|SONSTIGE HYPERPHENYLALANINAEMIEN
C2878662|T037|T43.692S|ICD10CM|POISONING BY OTHER PSYCHOSTIMULANTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH PSYCHOSTIMULANTS, SELF-HARM, SEQUELA
C2901902|T047|M86.549|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED HAND|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED HAND
C2901901|T047|M86.542|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, LEFT HAND|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, LEFT HAND
C2901900|T047|M86.541|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, RIGHT HAND|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, RIGHT HAND
C2887918|T047||ICD10CM|ALCOHOLIC HEPATIC FAILURE WITH COMA
C2887917|T047|K70.40|ICD10CM|ALCOHOLIC HEPATIC FAILURE WITHOUT COMA|ALCOHOLIC HEPATIC FAILURE WITHOUT COMA
C2854011|T191|C84.A9|ICD10CM|CUTANEOUS T-CELL LYMPHOMA, UNSPECIFIED, EXTRANODAL AND SOLID ORGAN SITES|CUTAN T-CELL LYMPHOMA, UNSP, EXTRNOD AND SOLID ORGAN SITES
C2854010|T191|C84.A8|ICD10CM|CUTANEOUS T-CELL LYMPHOMA, UNSPECIFIED, LYMPH NODES OF MULTIPLE SITES|CUTANEOUS T-CELL LYMPHOMA, UNSP, LYMPH NODES MULT SITE
C2869817|T037|S98.139S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF ONE UNSPECIFIED LESSER TOE, SEQUELA|COMPLETE TRAUMATIC AMP OF ONE UNSP LESSER TOE, SEQUELA
C2854003|T191|C84.A1|ICD10CM|CUTANEOUS T-CELL LYMPHOMA, UNSPECIFIED LYMPH NODES OF HEAD, FACE, AND NECK|CUTAN T-CELL LYMPHOMA, UNSP NODES OF HEAD, FACE, AND NECK
C2854002|T191|C84.A0|ICD10CM|CUTANEOUS T-CELL LYMPHOMA, UNSPECIFIED, UNSPECIFIED SITE|CUTANEOUS T-CELL LYMPHOMA, UNSPECIFIED, UNSPECIFIED SITE
C2854005|T191|C84.A3|ICD10CM|CUTANEOUS T-CELL LYMPHOMA, UNSPECIFIED, INTRA-ABDOMINAL LYMPH NODES|CUTANEOUS T-CELL LYMPHOMA, UNSP, INTRA-ABDOMINAL LYMPH NODES
C2854004|T191|C84.A2|ICD10CM|CUTANEOUS T-CELL LYMPHOMA, UNSPECIFIED, INTRATHORACIC LYMPH NODES|CUTANEOUS T-CELL LYMPHOMA, UNSP, INTRATHORACIC LYMPH NODES
C2854007|T191|C84.A5|ICD10CM|CUTANEOUS T-CELL LYMPHOMA, UNSPECIFIED, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|CUTAN T-CELL LYMPH, UNSP, NODES OF ING REGION AND LOWER LIMB
C2854006|T191|C84.A4|ICD10CM|CUTANEOUS T-CELL LYMPHOMA, UNSPECIFIED, LYMPH NODES OF AXILLA AND UPPER LIMB|CUTAN T-CELL LYMPHOMA, UNSP, NODES OF AXILLA AND UPPER LIMB
C2854009|T191|C84.A7|ICD10CM|CUTANEOUS T-CELL LYMPHOMA, UNSPECIFIED, SPLEEN|CUTANEOUS T-CELL LYMPHOMA, UNSPECIFIED, SPLEEN
C2854008|T191|C84.A6|ICD10CM|CUTANEOUS T-CELL LYMPHOMA, UNSPECIFIED, INTRAPELVIC LYMPH NODES|CUTANEOUS T-CELL LYMPHOMA, UNSP, INTRAPELVIC LYMPH NODES
C2869816|T037|S98.139D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF ONE UNSPECIFIED LESSER TOE, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF ONE UNSP LESSER TOE, SUBS
C2869815|T037|S98.139A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF ONE UNSPECIFIED LESSER TOE, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF ONE UNSP LESSER TOE, INIT
C2833182|T037|S12.040A|ICD10CM|DISPLACED LATERAL MASS FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED LATERAL MASS FX FIRST CERVCAL VERTEBRA, INIT
C2833183|T037|S12.040B|ICD10CM|DISPLACED LATERAL MASS FRACTURE OF FIRST CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISPL LATERAL MASS FX FIRST CERVCAL VERT, INIT FOR OPN FX
C2832519|T037|S06.6X2S|ICD10CM|TRAUMATIC SUBARACHNOID HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|TRAUM SUBRAC HEM W LOC OF 31-59 MIN, SEQUELA
C2886432|T037|T71.192S|ICD10CM|ASPHYXIATION DUE TO MECHANICAL THREAT TO BREATHING DUE TO OTHER CAUSES, INTENTIONAL SELF-HARM, SEQUELA|ASPHYX D/T MECH THRT TO BREATHE D/T OTH CAUSE, SLF-HRM, SQLA
C2902426|T047|M90.512|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, LEFT SHOULDER|OSTEONECROSIS IN DISEASES CLASSD ELSWHR, LEFT SHOULDER
C2902425|T047|M90.511|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, RIGHT SHOULDER|OSTEONECROSIS IN DISEASES CLASSD ELSWHR, RIGHT SHOULDER
C2902427|T047|M90.519|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, UNSPECIFIED SHOULDER|OSTEONECROSIS IN DISEASES CLASSD ELSWHR, UNSP SHOULDER
C2349331|T191|C7A.098|ICD10CM|MALIGNANT CARCINOID TUMORS OF OTHER SITES|MALIGNANT CARCINOID TUMORS OF OTHER SITES
C2886430|T037|T71.192A|ICD10CM|ASPHYXIATION DUE TO MECHANICAL THREAT TO BREATHING DUE TO OTHER CAUSES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|ASPHYX D/T MECH THRT TO BREATHE D/T OTH CAUSE, SLF-HRM, INIT
C2349326|T191|C7A.090|ICD10CM|MALIGNANT CARCINOID TUMOR OF THE BRONCHUS AND LUNG|MALIGNANT CARCINOID TUMOR OF THE BRONCHUS AND LUNG
C1336746|T191||ICD10CM|MALIGNANT CARCINOID TUMOR OF THE THYMUS
C2062573|T191||ICD10CM|MALIGNANT CARCINOID TUMOR OF THE STOMACH
C2349327|T191||ICD10CM|MALIGNANT CARCINOID TUMOR OF THE KIDNEY
C4270805|T191|C7A.094|ICD10CM|MALIGNANT CARCINOID TUMOR OF THE FOREGUT, UNSPECIFIED|MALIGNANT CARCINOID TUMOR OF THE FOREGUT, UNSPECIFIED
C4267837|T191|C7A.095|ICD10CM|MALIGNANT CARCINOID TUMOR OF THE MIDGUT, UNSPECIFIED|MALIGNANT CARCINOID TUMOR OF THE MIDGUT, UNSPECIFIED
C4267838|T191|C7A.096|ICD10CM|MALIGNANT CARCINOID TUMOR OF THE HINDGUT, UNSPECIFIED|MALIGNANT CARCINOID TUMOR OF THE HINDGUT, UNSPECIFIED
C2889601|T047|M08.812|ICD10CM|OTHER JUVENILE ARTHRITIS, LEFT SHOULDER|OTHER JUVENILE ARTHRITIS, LEFT SHOULDER
C2889600|T047|M08.811|ICD10CM|OTHER JUVENILE ARTHRITIS, RIGHT SHOULDER|OTHER JUVENILE ARTHRITIS, RIGHT SHOULDER
C2890567|T037|T84.093A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTERNAL LEFT KNEE PROSTHESIS, INITIAL ENCOUNTER|MECH COMPL OF INTERNAL LEFT KNEE PROSTHESIS, INIT ENCNTR
C2889602|T047|M08.819|ICD10CM|OTHER JUVENILE ARTHRITIS, UNSPECIFIED SHOULDER|OTHER JUVENILE ARTHRITIS, UNSPECIFIED SHOULDER
C2837912|T037|S32.411A|ICD10CM|DISPLACED FRACTURE OF ANTERIOR WALL OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF ANTERIOR WALL OF RIGHT ACETABULUM, INIT
C2837913|T037|S32.411B|ICD10CM|DISPLACED FRACTURE OF ANTERIOR WALL OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISP FX OF ANTERIOR WALL OF RIGHT ACETAB, INIT FOR OPN FX
C4268068|T047|E11.3211|ICD10CM|TYPE 2 DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, RIGHT EYE|TYPE 2 DIAB WITH MILD NONP RTNOP WITH MACULAR EDEMA, R EYE
C2874720|T048|F16.988|ICD10CM|HALLUCINOGEN USE, UNSPECIFIED WITH OTHER HALLUCINOGEN-INDUCED DISORDER|HALLUCINOGEN USE, UNSP W OTH HALLUCINOGEN-INDUCED DISORDER
C4268070|T047|E11.3213|ICD10CM|TYPE 2 DIABETES MELLITUS WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITH MACULAR EDEMA, BILATERAL|TYPE 2 DIABETES WITH MILD NONP RTNOP WITH MACULAR EDEMA, BI
C2500970|T060|B402|ICD10PCS|PULMONARY BLASTOMYCOSIS, UNSPECIFIED|IMAGING @ LOWER ARTERIES @ PLAIN RADIOGRAPHY @ HEPATIC ARTERY
C2832162|T037|S06.326S|ICD10CM|CONTUSION AND LACERATION OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|CONTUS/LAC L CEREB W LOC >24 HR W/O RET CONSC W SURV, SQLA
C2500963|T060|B400|ICD10PCS|ACUTE PULMONARY BLASTOMYCOSIS|IMAGING @ LOWER ARTERIES @ PLAIN RADIOGRAPHY @ ABDOMINAL AORTA
C0343920|T047|B40.1|DMDICD10|CHRONIC PULMONARY BLASTOMYCOSIS|CHRONISCHE BLASTOMYKOSE DER LUNGE
C2874719|T048|F16.983|ICD10CM|HALLUCINOGEN USE, UNSPECIFIED WITH HALLUCINOGEN PERSISTING PERCEPTION DISORDER (FLASHBACKS)|HALLUCIGN USE, UNSP W HALLUCIGN PERSIST PERCEPTION DISORDER
C4237363|T048|F16.980|ICD10CM|HALLUCINOGEN USE, UNSPECIFIED WITH HALLUCINOGEN-INDUCED ANXIETY DISORDER|PHENCYCLIDINE INDUCED ANXIETY DISORDER, WITHOUT USE DISORDER
C0840000|T047|M86.8X2|ICD10CM|OTHER OSTEOMYELITIS, UPPER ARM|OTHER OSTEOMYELITIS, UPPER ARM
C2889373|T047|M05.851|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT HIP|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT HIP
C2889374|T047|M05.852|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HIP|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HIP
C2901933|T047|M86.8X1|ICD10CM|OTHER OSTEOMYELITIS, SHOULDER|OTHER OSTEOMYELITIS, SHOULDER
C2889375|T047|M05.859|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED HIP|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSP HIP
C0839998|T047|M86.8X0|ICD10CM|OTHER OSTEOMYELITIS, MULTIPLE SITES|OTHER OSTEOMYELITIS, MULTIPLE SITES
C2901437|T046|M84.634A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, LEFT RADIUS, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE IN OTH DISEASE, LEFT RADIUS, INIT
C2832633|T037|S06.890S|ICD10CM|OTHER SPECIFIED INTRACRANIAL INJURY WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|OTH INTRACRANIAL INJURY W/O LOSS OF CONSCIOUSNESS, SEQUELA
C2837810|T037|S32.302A|ICD10CM|UNSPECIFIED FRACTURE OF LEFT ILIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF LEFT ILIUM, INIT ENCNTR FOR CLOSED FRACTURE
C2837811|T037|S32.302B|ICD10CM|UNSPECIFIED FRACTURE OF LEFT ILIUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF LEFT ILIUM, INIT ENCNTR FOR OPEN FRACTURE
C2896514|T046|M80.022A|ICD10CM|AGE-RELATED OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, LEFT HUMERUS, INITIAL ENCOUNTER FOR FRACTURE|AGE-REL OSTEOPOR W CURRENT PATH FRACTURE, L HUMERUS, INIT
C2889162|T047|M05.172|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT|RHEU LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT ANK/FT
C2832631|T037|S06.890A|ICD10CM|OTHER SPECIFIED INTRACRANIAL INJURY WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|INTCRAN INJ W/O LOSS OF CONSCIOUSNESS, INIT ENCNTR
C2882728|T047|I70.245|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF LEFT LEG WITH ULCERATION OF OTHER PART OF FOOT|ATHSCL NATIVE ARTERIES OF LEFT LEG W ULCERATION OTH PRT FOOT
C0349337|T048||ICD10CM|OTHER PHOBIC ANXIETY DISORDERS
C0349231|T048|F40|DMDICD10|PHOBIC ANXIETY DISORDER, UNSPECIFIED|PHOBISCHE STOERUNGEN
C2830359|T033|R40.2124|ICD10CM|COMA SCALE, EYES OPEN, TO PAIN, 24 HOURS OR MORE AFTER HOSPITAL ADMISSION|COMA SCALE, EYES OPEN, TO PAIN, 24+HRS
C2889161|T047|M05.171|ICD10CM|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT|RHEU LUNG DISEASE W RHEUMATOID ARTHRITIS OF RIGHT ANK/FT
C2856999|T037|S72.064A|ICD10CM|NONDISPLACED ARTICULAR FRACTURE OF HEAD OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISPLACED ARTICULAR FRACTURE OF HEAD OF RIGHT FEMUR, INIT
C2857001|T037|S72.064C|ICD10CM|NONDISPLACED ARTICULAR FRACTURE OF HEAD OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP ARTIC FX HEAD OF R FEMR, INIT FOR OPN FX TYPE 3A/B/C
C2857000|T037|S72.064B|ICD10CM|NONDISPLACED ARTICULAR FRACTURE OF HEAD OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP ARTIC FX HEAD OF R FEMUR, INIT FOR OPN FX TYPE I/2
C2830355|T033|R40.2120|ICD10CM|COMA SCALE, EYES OPEN, TO PAIN, UNSPECIFIED TIME|COMA SCALE, EYES OPEN, TO PAIN, UNSPECIFIED TIME
C2830356|T033|R40.2121|ICD10CM|COMA SCALE, EYES OPEN, TO PAIN, IN THE FIELD [EMT OR AMBULANCE]|COMA SCALE, EYES OPEN, TO PAIN, IN THE FIELD
C2830357|T033|R40.2122|ICD10CM|COMA SCALE, EYES OPEN, TO PAIN, AT ARRIVAL TO EMERGENCY DEPARTMENT|COMA SCALE, EYES OPEN, TO PAIN, EMR
C0840019|T037|M87.19|ICD10CM|OSTEONECROSIS DUE TO DRUGS, MULTIPLE SITES|OSTEONECROSIS DUE TO DRUGS, MULTIPLE SITES
C2855935|T037|S68.127S|ICD10CM|PARTIAL TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF LEFT LITTLE FINGER, SEQUELA|PARTIAL TRAUMATIC MCP AMPUTATION OF L LITTLE FINGER, SEQUELA
C2830358|T033|R40.2123|ICD10CM|COMA SCALE, EYES OPEN, TO PAIN, AT HOSPITAL ADMISSION|COMA SCALE, EYES OPEN, TO PAIN, AT HOSPITAL ADMISSION
C2882792|T047|I70.363|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, BILATERAL LEGS|ATHSCL UNSP TYPE BYPASS OF THE EXTRM W GANGRENE, BI LEGS
C2882791|T047|I70.362|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, LEFT LEG|ATHSCL UNSP TYPE BYPASS OF THE EXTRM W GANGRENE, LEFT LEG
C2882790|T047|I70.361|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, RIGHT LEG|ATHSCL UNSP TYPE BYPASS OF THE EXTRM W GANGRENE, RIGHT LEG
C2889193|T047|M05.272|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF LEFT ANK/FT
C2889194|T047|M05.279|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF UNSP ANK/FT
C2882794|T047|I70.369|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, UNSPECIFIED EXTREMITY|ATHSCL UNSP TYPE BYPASS OF THE EXTRM W GANGRENE, UNSP EXTRM
C2882793|T047|I70.368|ICD10CM|ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES WITH GANGRENE, OTHER EXTREMITY|ATHSCL UNSP TYPE BYPASS OF THE EXTRM W GANGRENE, OTH EXTRM
C2901985|T046|M87.10|ICD10CM|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED BONE|OSTEONECROSIS DUE TO DRUGS, UNSPECIFIED BONE
C4270212|T046|T83.028A|ICD10CM|DISPLACEMENT OF OTHER URINARY CATHETER, INITIAL ENCOUNTER|DISPLACEMENT OF OTHER URINARY CATHETER, INITIAL ENCOUNTER
C2835377|T037|S22.061A|ICD10CM|STABLE BURST FRACTURE OF T7-T8 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|STABLE BURST FRACTURE OF T7-T8 VERTEBRA, INIT FOR CLOS FX
C2857753|T037|S72.323A|ICD10CM|DISPLACED TRANSVERSE FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED TRANSVERSE FRACTURE OF SHAFT OF UNSP FEMUR, INIT
C2857755|T037|S72.323C|ICD10CM|DISPLACED TRANSVERSE FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL TRANSVERSE FX SHAFT OF UNSP FEMR, 7THC
C2857754|T037|S72.323B|ICD10CM|DISPLACED TRANSVERSE FRACTURE OF SHAFT OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPL TRANSVERSE FX SHAFT OF UNSP FEMR, 7THB
C2887838|T047|K51.90|ICD10CM|ULCERATIVE COLITIS, UNSPECIFIED, WITHOUT COMPLICATIONS|ULCERATIVE COLITIS, UNSPECIFIED, WITHOUT COMPLICATIONS
C2874557|T048|F13.930|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH WITHDRAWAL, UNCOMPLICATED|SEDATV/HYP/ANXIOLYTC USE, UNSP W WITHDRAWAL, UNCOMPLICATED
C2874558|T048|F13.931|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH WITHDRAWAL DELIRIUM|SEDATV/HYP/ANXIOLYTC USE, UNSP W WITHDRAWAL DELIRIUM
C2874559|T048|F13.932|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH WITHDRAWAL WITH PERCEPTUAL DISTURBANCES|SEDATV/HYP/ANXIOLYTC USE, UNSP W W/DRAWAL W PERCEPTL DISTURB
C2874560|T048|F13.939|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH WITHDRAWAL, UNSPECIFIED|SEDATV/HYP/ANXIOLYTC USE, UNSP W WITHDRAWAL, UNSP
C0348353|T191|C45.7|DMDICD10|MESOTHELIOMA OF OTHER SITES|MESOTHELIOM SONSTIGER LOKALISATIONEN
C2838675|T037|S34.123D|ICD10CM|INCOMPLETE LESION OF L3 LEVEL OF LUMBAR SPINAL CORD, SUBSEQUENT ENCOUNTER|INCOMPLETE LESION OF L3 LEVEL OF LUMBAR SPINAL CORD, SUBS
C2838674|T037|S34.123A|ICD10CM|INCOMPLETE LESION OF L3 LEVEL OF LUMBAR SPINAL CORD, INITIAL ENCOUNTER|INCOMPLETE LESION OF L3 LEVEL OF LUMBAR SPINAL CORD, INIT
C2837568|T037|S32.032B|ICD10CM|UNSTABLE BURST FRACTURE OF THIRD LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSTABLE BURST FX THIRD LUM VERTEBRA, INIT FOR OPN FX
C2901538|T046|M84.669A|ICD10CM|PATHOLOGICAL FRACTURE IN OTHER DISEASE, UNSPECIFIED TIBIA AND FIBULA, INITIAL ENCOUNTER FOR FRACTURE|PATH FRACTURE IN OTH DISEASE, UNSP TIBIA AND FIBULA, INIT
C2838676|T037|S34.123S|ICD10CM|INCOMPLETE LESION OF L3 LEVEL OF LUMBAR SPINAL CORD, SEQUELA|INCOMPLETE LESION OF L3 LEVEL OF LUMBAR SPINAL CORD, SEQUELA
C0600327|T047|A48.3|DMDICD10|TOXIC SHOCK SYNDROME|SYNDROM DES TOXISCHEN SCHOCKS
C0023241|T047|A48.1|DMDICD10|LEGIONNAIRES' DISEASE|LEGIONELLOSE MIT PNEUMONIE
C2887103|T047|A48.0|ICD10CM|GAS GANGRENE|CLOSTRIDIAL CELLULITIS
C2845894|T191|C65.9|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED RENAL PELVIS|MALIGNANT NEOPLASM OF UNSPECIFIED RENAL PELVIS
C2832511|T037|S06.6X0S|ICD10CM|TRAUMATIC SUBARACHNOID HEMORRHAGE WITHOUT LOSS OF CONSCIOUSNESS, SEQUELA|TRAUM SUBRAC HEM W/O LOSS OF CONSCIOUSNESS, SEQUELA
C2885221|T037|T62.0X2A|ICD10CM|TOXIC EFFECT OF INGESTED MUSHROOMS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF INGESTED MUSHROOMS, SELF-HARM, INIT
C2845893|T191|C65.1|ICD10CM|MALIGNANT NEOPLASM OF RIGHT RENAL PELVIS|MALIGNANT NEOPLASM OF RIGHT RENAL PELVIS
C0864886|T191|C30.0|ICD10CM|MALIGNANT NEOPLASM OF NASAL CAVITY|MALIGNANT NEOPLASM OF INTERNAL NOSE
C2837942|T191|C30.1|ICD10CM|MALIGNANT NEOPLASM OF MIDDLE EAR|MALIGNANT NEOPLASM OF INNER EAR
C2832509|T037|S06.6X0A|ICD10CM|TRAUMATIC SUBARACHNOID HEMORRHAGE WITHOUT LOSS OF CONSCIOUSNESS, INITIAL ENCOUNTER|TRAUM SUBRAC HEM W/O LOSS OF CONSCIOUSNESS, INIT
C3264001|T047|G40.B11|ICD10CM|JUVENILE MYOCLONIC EPILEPSY, INTRACTABLE, WITH STATUS EPILEPTICUS|JUVENILE MYOCLONIC EPILEPSY, INTRACTABLE, W STAT EPI
C2843308|T037|S48.121A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEVEL BETWEEN RIGHT SHOULDER AND ELBOW, INITIAL ENCOUNTER|PARTIAL TRAUM AMP AT LEVEL BETW R SHOULDER AND ELBOW, INIT
C2859096|T037|S72.91XA|ICD10CM|UNSPECIFIED FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF RIGHT FEMUR, INIT FOR CLOS FX
C2859098|T037|S72.91XC|ICD10CM|UNSPECIFIED FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP FRACTURE OF RIGHT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C3264002|T047|G40.B19|ICD10CM|JUVENILE MYOCLONIC EPILEPSY, INTRACTABLE, WITHOUT STATUS EPILEPTICUS|JUVENILE MYOCLONIC EPILEPSY, INTRACTABLE, W/O STAT EPI
C2856057|T037|S68.623S|ICD10CM|PARTIAL TRAUMATIC TRANSPHALANGEAL AMPUTATION OF LEFT MIDDLE FINGER, SEQUELA|PARTIAL TRAUMATIC TRNSPHAL AMP OF L MID FINGER, SEQUELA
C3887878|T047|E06.5|ICD10CM|OTHER CHRONIC THYROIDITIS|CHRONIC FIBROUS THYROIDITIS
C0342179|T046|E06.4|DMDICD10|DRUG-INDUCED THYROIDITIS|ARZNEIMITTELINDUZIERTE THYREOIDITIS
C1406948|T047||ICD10CM|SUBACUTE THYROIDITIS
C0494612|T020|I66.9|DMDICD10|OCCLUSION AND STENOSIS OF UNSPECIFIED CEREBRAL ARTERY|VERSCHLUSS UND STENOSE NICHT NAEHER BEZEICHNETER INTRAKRANIELLER ARTERIE
C0920350|T047|E06.3|DMDICD10|AUTOIMMUNE THYROIDITIS|AUTOIMMUNTHYREOIDITIS
C0342178|T047|E06.2|DMDICD10|CHRONIC THYROIDITIS WITH TRANSIENT THYROTOXICOSIS|CHRONISCHE THYREOIDITIS MIT TRANSITORISCHER HYPERTHYREOSE
C0040147|T047|E06.9|DMDICD10|THYROIDITIS, UNSPECIFIED|THYREOIDITIS, NICHT NAEHER BEZEICHNET
C2858870|T037|S72.462C|ICD10CM|DISPLACED SUPRACONDYLAR FRACTURE WITH INTRACONDYLAR EXTENSION OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPL SUPRCNDL FX W INTRCNDL EXTN LOW END L FEMR, 7THC
C2889894|T037|T82.310A|ICD10CM|BREAKDOWN (MECHANICAL) OF AORTIC (BIFURCATION) GRAFT (REPLACEMENT), INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF AORTIC (BIFURCATION) GRAFT, INIT
C2875345|T047|G83.12|ICD10CM|MONOPLEGIA OF LOWER LIMB AFFECTING LEFT DOMINANT SIDE|MONOPLEGIA OF LOWER LIMB AFFECTING LEFT DOMINANT SIDE
C2874640|T048|F15.182|ICD10CM|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED SLEEP DISORDER|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED SLEEP DISORDER
C0375224|T184|G83.10|ICD10CM|MONOPLEGIA OF LOWER LIMB AFFECTING UNSPECIFIED SIDE|MONOPLEGIA OF LOWER LIMB AFFECTING UNSPECIFIED SIDE
C2874638|T048|F15.180|ICD10CM|OTHER STIMULANT ABUSE WITH STIMULANT-INDUCED ANXIETY DISORDER|OTH STIMULANT ABUSE WITH STIMULANT-INDUCED ANXIETY DISORDER
C2875347|T047|G83.14|ICD10CM|MONOPLEGIA OF LOWER LIMB AFFECTING LEFT NONDOMINANT SIDE|MONOPLEGIA OF LOWER LIMB AFFECTING LEFT NONDOMINANT SIDE
C4268247|T048|F15.188|ICD10CM|OTHER STIMULANT ABUSE WITH OTHER STIMULANT-INDUCED DISORDER|AMPHETAMINE OR OTHER STIMULANT USE DISORDER, MILD, WITH AMPHETAMINE OR OTHER STIMULANT INDUCED OBSESSIVE-COMPULSIVE OR RELATED DISORDER
C3263971|T047|G40.509|ICD10CM|EPILEPTIC SEIZURES RELATED TO EXTERNAL CAUSES, NOT INTRACTABLE, WITHOUT STATUS EPILEPTICUS|EPILEPTIC SEIZ REL TO EXTRN CAUSES, NOT NTRCT, W/O STAT EPI
C4268788|T046|M84.756A|ICD10CM|COMPLETE TRANSVERSE ATYPICAL FEMORAL FRACTURE, UNSPECIFIED LEG, INITIAL ENCOUNTER FOR FRACTURE|COMPLETE TRANSVERSE ATYP FEMORAL FRACTURE, UNSP LEG, INIT
C3263969|T047|G40.501|ICD10CM|EPILEPTIC SEIZURES RELATED TO EXTERNAL CAUSES, NOT INTRACTABLE, WITH STATUS EPILEPTICUS|EPILEPTIC SEIZ REL TO EXTRN CAUSES, NOT NTRCT, W STAT EPI
C0152946|T047|A22.7|DMDICD10|ANTHRAX SEPSIS|MILZBRANDSEPSIS
C1411077|T047||ICD10CM|PULMONARY ANTHRAX
C0686396|T191|C79.32|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF CEREBRAL MENINGES|SECONDARY MALIGNANT NEOPLASM OF CEREBRAL MENINGES
C0220650|T191|C79.31|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF BRAIN|SECONDARY MALIGNANT NEOPLASM OF BRAIN
C2886137|T037|T65.812S|ICD10CM|TOXIC EFFECT OF LATEX, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF LATEX, INTENTIONAL SELF-HARM, SEQUELA
C2842043|T191|C49.10|ICD10CM|MALIGNANT NEOPLASM OF CONNECTIVE AND SOFT TISSUE OF UNSPECIFIED UPPER LIMB, INCLUDING SHOULDER|MALIG NEOPLM OF CONN & SOFT TISS OF UNSP UPR LMB, INC SHLDR
C2842044|T191|C49.11|ICD10CM|MALIGNANT NEOPLASM OF CONNECTIVE AND SOFT TISSUE OF RIGHT UPPER LIMB, INCLUDING SHOULDER|MALIG NEOPLM OF CONN AND SOFT TISS OF R UPR LIMB, INC SHLDR
C2842045|T191|C49.12|ICD10CM|MALIGNANT NEOPLASM OF CONNECTIVE AND SOFT TISSUE OF LEFT UPPER LIMB, INCLUDING SHOULDER|MALIG NEOPLM OF CONN AND SOFT TISS OF L UPR LIMB, INC SHLDR
C2886135|T037|T65.812A|ICD10CM|TOXIC EFFECT OF LATEX, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF LATEX, INTENTIONAL SELF-HARM, INIT ENCNTR
C2853857|T191|C82.68|ICD10CM|CUTANEOUS FOLLICLE CENTER LYMPHOMA, LYMPH NODES OF MULTIPLE SITES|CUTANEOUS FOLLICLE CENTER LYMPHOMA, LYMPH NODES MULT SITE
C3647898|T191|C82.69|ICD10CM|CUTANEOUS FOLLICLE CENTER LYMPHOMA, EXTRANODAL AND SOLID ORGAN SITES|CUTAN FOLICL CENTER LYMPHOMA, EXTRNOD AND SOLID ORGAN SITES
C0477394|T047|G62.8|ICD10CM|OTHER SPECIFIED POLYNEUROPATHIES|OTHER SPECIFIED POLYNEUROPATHIES
C3648008|T191|C82.62|ICD10CM|CUTANEOUS FOLLICLE CENTER LYMPHOMA, INTRATHORACIC LYMPH NODES|CUTANEOUS FOLLICLE CENTER LYMPHOMA, INTRATHORAC LYMPH NODES
C3648010|T191|C82.63|ICD10CM|CUTANEOUS FOLLICLE CENTER LYMPHOMA, INTRA-ABDOMINAL LYMPH NODES|CUTANEOUS FOLLICLE CENTER LYMPHOMA, INTRA-ABD LYMPH NODES
C2853849|T191|C82.60|ICD10CM|CUTANEOUS FOLLICLE CENTER LYMPHOMA, UNSPECIFIED SITE|CUTANEOUS FOLLICLE CENTER LYMPHOMA, UNSPECIFIED SITE
C3648011|T191|C82.61|ICD10CM|CUTANEOUS FOLLICLE CENTER LYMPHOMA, LYMPH NODES OF HEAD, FACE, AND NECK|CUTAN FOLICL CENTER LYMPHOMA, NODES OF HEAD, FACE, AND NECK
C2875306|T047||ICD10CM|RADIATION-INDUCED POLYNEUROPATHY
C2853856|T191|C82.67|ICD10CM|CUTANEOUS FOLLICLE CENTER LYMPHOMA, SPLEEN|CUTANEOUS FOLLICLE CENTER LYMPHOMA, SPLEEN
C3648034|T191|C82.64|ICD10CM|CUTANEOUS FOLLICLE CENTER LYMPHOMA, LYMPH NODES OF AXILLA AND UPPER LIMB|CUTAN FOLICL CENTER LYMPHOMA, NODES OF AXILLA AND UPPER LIMB
C1135343|T047|G62.81|ICD10CM|CRITICAL ILLNESS POLYNEUROPATHY|ACUTE MOTOR NEUROPATHY
C2860186|T037|S79.131A|ICD10CM|SALTER-HARRIS TYPE III PHYSEAL FRACTURE OF LOWER END OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|SLTR-HARIS TYPE III PHYSEAL FX LOWER END OF R FEMUR, INIT
C2869830|T037|S98.149S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF ONE UNSPECIFIED LESSER TOE, SEQUELA|PARTIAL TRAUMATIC AMPUTATION OF ONE UNSP LESSER TOE, SEQUELA
C2859994|T037|S78.029S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT UNSPECIFIED HIP JOINT, SEQUELA|PARTIAL TRAUMATIC AMPUTATION AT UNSP HIP JOINT, SEQUELA
C2887826|T047|K51.513|ICD10CM|LEFT SIDED COLITIS WITH FISTULA|LEFT SIDED COLITIS WITH FISTULA
C2887825|T047|K51.512|ICD10CM|LEFT SIDED COLITIS WITH INTESTINAL OBSTRUCTION|LEFT SIDED COLITIS WITH INTESTINAL OBSTRUCTION
C2887824|T047|K51.511|ICD10CM|LEFT SIDED COLITIS WITH RECTAL BLEEDING|LEFT SIDED COLITIS WITH RECTAL BLEEDING
C2887827|T047|K51.514|ICD10CM|LEFT SIDED COLITIS WITH ABSCESS|LEFT SIDED COLITIS WITH ABSCESS
C2887829|T047|K51.519|ICD10CM|LEFT SIDED COLITIS WITH UNSPECIFIED COMPLICATIONS|LEFT SIDED COLITIS WITH UNSPECIFIED COMPLICATIONS
C2887828|T047|K51.518|ICD10CM|LEFT SIDED COLITIS WITH OTHER COMPLICATION|LEFT SIDED COLITIS WITH OTHER COMPLICATION
C2874864|T048||ICD10CM|MANIC EPISODE WITHOUT PSYCHOTIC SYMPTOMS, MILD
C2874863|T048|F30.10|ICD10CM|MANIC EPISODE WITHOUT PSYCHOTIC SYMPTOMS, UNSPECIFIED|MANIC EPISODE WITHOUT PSYCHOTIC SYMPTOMS, UNSPECIFIED
C2874866|T048||ICD10CM|MANIC EPISODE, SEVERE, WITHOUT PSYCHOTIC SYMPTOMS
C2874865|T048||ICD10CM|MANIC EPISODE WITHOUT PSYCHOTIC SYMPTOMS, MODERATE
C2832242|T037|S06.345S|ICD10CM|TRAUMATIC HEMORRHAGE OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, SEQUELA|TRAUM HEMOR R CEREB W LOC >24 HR W RET CONSC LEV, SEQUELA
C2889935|T037|T82.330A|ICD10CM|LEAKAGE OF AORTIC (BIFURCATION) GRAFT (REPLACEMENT), INITIAL ENCOUNTER|LEAKAGE OF AORTIC (BIFURCATION) GRAFT (REPLACEMENT), INIT
C4267945|T047|E08.3591|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH PROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|DIAB WITH PROLIF DIABETIC RTNOP WITHOUT MACULAR EDEMA, R EYE
C2885107|T037|T60.92XA|ICD10CM|TOXIC EFFECT OF UNSPECIFIED PESTICIDE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF UNSP PESTICIDE, INTENTIONAL SELF-HARM, INIT
C2838101|T037|S32.432B|ICD10CM|DISPLACED FRACTURE OF ANTERIOR COLUMN [ILIOPUBIC] OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|DISP FX OF ANTERIOR COLUMN OF LEFT ACETAB, INIT FOR OPN FX
C2838100|T037|S32.432A|ICD10CM|DISPLACED FRACTURE OF ANTERIOR COLUMN [ILIOPUBIC] OF LEFT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF ANTERIOR COLUMN OF LEFT ACETABULUM, INIT
C4268383|T047|H35.3222|ICD10CM|EXUDATIVE AGE-RELATED MACULAR DEGENERATION, LEFT EYE, WITH INACTIVE CHOROIDAL NEOVASCULARIZATION|EXDTVE AGE-REL MCLR DEGN, LEFT EYE, WITH INACT CHRDL NEOVAS
C4268384|T047|H35.3223|ICD10CM|EXUDATIVE AGE-RELATED MACULAR DEGENERATION, LEFT EYE, WITH INACTIVE SCAR|EXUDATIVE AGE-REL MCLR DEGN, LEFT EYE, WITH INACTIVE SCAR
C4268381|T047|H35.3220|ICD10CM|EXUDATIVE AGE-RELATED MACULAR DEGENERATION, LEFT EYE, STAGE UNSPECIFIED|EXUDATIVE AGE-RELATED MCLR DEGN, LEFT EYE, STAGE UNSPECIFIED
C4268382|T047|H35.3221|ICD10CM|EXUDATIVE AGE-RELATED MACULAR DEGENERATION, LEFT EYE, WITH ACTIVE CHOROIDAL NEOVASCULARIZATION|EXDTVE AGE-REL MCLR DEGN, LEFT EYE, WITH ACTV CHRDL NEOVAS
C2885109|T037|T60.92XS|ICD10CM|TOXIC EFFECT OF UNSPECIFIED PESTICIDE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF UNSP PESTICIDE, SELF-HARM, SEQUELA
C0041948|T047||ICD10CM|UNSPECIFIED KIDNEY FAILURE
C2882105|T047|I21.19|ICD10CM|ST ELEVATION (STEMI) MYOCARDIAL INFARCTION INVOLVING OTHER CORONARY ARTERY OF INFERIOR WALL|STEMI INVOLVING OTH CORONARY ARTERY OF INFERIOR WALL
C2882557|T047|I69.269|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING UNSPECIFIED SIDE|OTH PARLYT SYNDROME FOL OTH NTRM INTCRN HEMOR AFF UNSP SIDE
C2882555|T047|I69.264|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING LEFT NON-DOMINANT SIDE|OTH PARLYT SYND FOL OTH NTRM INTCRN HEMOR AFF L NONDOM SIDE
C2882556|T047|I69.265|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE, BILATERAL|OTH PARALYTIC SYNDROME FOLLOWING OTH NTRM INTCRN HEMOR, BI
C2882552|T047|I69.261|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING RIGHT DOMINANT SIDE|OTH PARLYT SYND FOL OTH NTRM INTCRN HEMOR AFF RIGHT DOM SIDE
C2882553|T047|I69.262|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING LEFT DOMINANT SIDE|OTH PARLYT SYND FOL OTH NTRM INTCRN HEMOR AFF LEFT DOM SIDE
C2882554|T047|I69.263|ICD10CM|OTHER PARALYTIC SYNDROME FOLLOWING OTHER NONTRAUMATIC INTRACRANIAL HEMORRHAGE AFFECTING RIGHT NON-DOMINANT SIDE|OTH PARLYT SYND FOL OTH NTRM INTCRN HEMOR AFF R NONDOM SIDE
C2876946|T037|T37.8X2S|ICD10CM|POISONING BY OTHER SPECIFIED SYSTEMIC ANTI-INFECTIVES AND ANTIPARASITICS, INTENTIONAL SELF-HARM, SEQUELA|POISN BY OTH SYSTEMIC ANTI-INFECT/PARASIT, SLF-HRM, SEQUELA
C0432482|T019|Q99.2|DMDICD10|FRAGILE X CHROMOSOME|FRAGILES X-CHROMOSOM
C2854096|T191||ICD10CM|PROLYMPHOCYTIC LEUKEMIA OF B-CELL TYPE, IN REMISSION
C2854095|T191|C91.30|ICD10CM|PROLYMPHOCYTIC LEUKEMIA OF B-CELL TYPE NOT HAVING ACHIEVED REMISSION|PROLYMPHOCYTIC LEUKEMIA OF B-CELL TYPE NOT ACHIEVE REMISSION
C2854097|T191||ICD10CM|PROLYMPHOCYTIC LEUKEMIA OF B-CELL TYPE, IN RELAPSE
C4270539|T046|T85.625A|ICD10CM|DISPLACEMENT OF OTHER NERVOUS SYSTEM DEVICE, IMPLANT OR GRAFT, INITIAL ENCOUNTER|DISPLACMNT OF NERVOUS SYS DEVICE, IMPLANT OR GRAFT, INIT
C0029816|T047|G70.89|ICD10CM|OTHER SPECIFIED MYONEURAL DISORDERS|OTHER SPECIFIED MYONEURAL DISORDERS
C2888840|T047|M00.139|ICD10CM|PNEUMOCOCCAL ARTHRITIS, UNSPECIFIED WRIST|PNEUMOCOCCAL ARTHRITIS, UNSPECIFIED WRIST
C2832667|T037|S06.899A|ICD10CM|OTHER SPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, INITIAL ENCOUNTER|INTCRAN INJ W LOSS OF CONSCIOUSNESS OF UNSP DURATION, INIT
C3250442|T047||ICD10CM|LAMBERT-EATON SYNDROME IN DISEASE CLASSIFIED ELSEWHERE
C3161080|T047|G70.80|ICD10CM|LAMBERT-EATON SYNDROME, UNSPECIFIED|LAMBERT-EATON SYNDROME, UNSPECIFIED
C2888838|T047|M00.131|ICD10CM|PNEUMOCOCCAL ARTHRITIS, RIGHT WRIST|PNEUMOCOCCAL ARTHRITIS, RIGHT WRIST
C2888839|T047|M00.132|ICD10CM|PNEUMOCOCCAL ARTHRITIS, LEFT WRIST|PNEUMOCOCCAL ARTHRITIS, LEFT WRIST
C2832160|T037|S06.326A|ICD10CM|CONTUSION AND LACERATION OF LEFT CEREBRUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|CONTUS/LAC L CEREB W LOC >24 HR W/O RET CONSC W SURV, INIT
C0477543|T047||ICD10CM|OTHER PSORIATIC ARTHROPATHY
C2889985|T037|T82.42XS|ICD10CM|DISPLACEMENT OF VASCULAR DIALYSIS CATHETER, SEQUELA|DISPLACEMENT OF VASCULAR DIALYSIS CATHETER, SEQUELA
C2888178|T047|L40.52|ICD10CM|PSORIATIC ARTHRITIS MUTILANS|PSORIATIC ARTHRITIS MUTILANS
C0343176|T047|L40.53|ICD10CM|PSORIATIC SPONDYLITIS|PSORIATIC SPONDYLITIS
C0003872|T047|L40.50|ICD10CM|ARTHROPATHIC PSORIASIS, UNSPECIFIED|ARTHROPATHIC PSORIASIS, UNSPECIFIED
C0409682|T047|L40.51|ICD10CM|DISTAL INTERPHALANGEAL PSORIATIC ARTHROPATHY|DISTAL INTERPHALANGEAL PSORIATIC ARTHROPATHY
C2888179|T047|L40.54|ICD10CM|PSORIATIC JUVENILE ARTHROPATHY|PSORIATIC JUVENILE ARTHROPATHY
C2889984|T037|T82.42XD|ICD10CM|DISPLACEMENT OF VASCULAR DIALYSIS CATHETER, SUBSEQUENT ENCOUNTER|DISPLACEMENT OF VASCULAR DIALYSIS CATHETER, SUBS ENCNTR
C2856655|T037|S72.025B|ICD10CM|NONDISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|NONDISP FX OF EPIPHY (SEPARATION) (UPPER) OF L FEMR, 7THB
C2856656|T037|S72.025C|ICD10CM|NONDISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP FX OF EPIPHY (SEPARATION) (UPPER) OF L FEMR, 7THC
C2889983|T037|T82.42XA|ICD10CM|DISPLACEMENT OF VASCULAR DIALYSIS CATHETER, INITIAL ENCOUNTER|DISPLACEMENT OF VASCULAR DIALYSIS CATHETER, INIT ENCNTR
C2856654|T037|S72.025A|ICD10CM|NONDISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF EPIPHY (SEPARATION) (UPPER) OF L FEMUR, INIT
C2885426|T037|T63.082S|ICD10CM|TOXIC EFFECT OF VENOM OF OTHER AFRICAN AND ASIAN SNAKE, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFF OF VENOM OF AFRICAN AND ASIAN SNAKE, SLF-HRM, SQLA
C2890879|T037|T84.625A|ICD10CM|INFECTION AND INFLAMMATORY REACTION DUE TO INTERNAL FIXATION DEVICE OF LEFT FIBULA, INITIAL ENCOUNTER|INFECT/INFLM REACTION DUE TO INT FIX OF LEFT FIBULA, INIT
C2910922|T033|Z48.290|ICD10CM|ENCOUNTER FOR AFTERCARE FOLLOWING BONE MARROW TRANSPLANT|ENCOUNTER FOR AFTERCARE FOLLOWING BONE MARROW TRANSPLANT
C2901863|T047|M86.371|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, RIGHT ANKLE AND FOOT|CHRONIC MULTIFOCAL OSTEOMYELITIS, RIGHT ANKLE AND FOOT
C2905771|T037|X79.XXXS|ICD10CM|INTENTIONAL SELF-HARM BY BLUNT OBJECT, SEQUELA|INTENTIONAL SELF-HARM BY BLUNT OBJECT, SEQUELA
C2901864|T047|M86.372|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, LEFT ANKLE AND FOOT|CHRONIC MULTIFOCAL OSTEOMYELITIS, LEFT ANKLE AND FOOT
C2901865|T047|M86.379|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, UNSPECIFIED ANKLE AND FOOT|CHRONIC MULTIFOCAL OSTEOMYELITIS, UNSPECIFIED ANKLE AND FOOT
C2838043|T037|S32.416B|ICD10CM|NONDISPLACED FRACTURE OF ANTERIOR WALL OF UNSPECIFIED ACETABULUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|NONDISP FX OF ANTERIOR WALL OF UNSP ACETAB, INIT FOR OPN FX
C2882622|T047|I69.841|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING RIGHT DOMINANT SIDE|MONOPLG LOW LMB FOL OTH CEREBVASC DISEASE AFF RIGHT DOM SIDE
C2882623|T047|I69.842|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING LEFT DOMINANT SIDE|MONOPLG LOW LMB FOL OTH CEREBVASC DISEASE AFF LEFT DOM SIDE
C2882624|T047|I69.843|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING RIGHT NON-DOMINANT SIDE|MONOPLG LOW LMB FOL OTH CEREBVASC DIS AFF RIGHT NONDOM SIDE
C2882625|T047|I69.844|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING LEFT NON-DOMINANT SIDE|MONOPLG LOW LMB FOL OTH CEREBVASC DIS AFF LEFT NONDOM SIDE
C2882626|T047|I69.849|ICD10CM|MONOPLEGIA OF LOWER LIMB FOLLOWING OTHER CEREBROVASCULAR DISEASE AFFECTING UNSPECIFIED SIDE|MONOPLG LOW LMB FOL OTH CEREBVASC DISEASE AFF UNSP SIDE
C2832507|T037|S06.5X9S|ICD10CM|TRAUMATIC SUBDURAL HEMORRHAGE WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|TRAUM SUBDR HEM W LOC OF UNSP DURATION, SEQUELA
C0153025|T047|B02.23|ICD10CM|POSTHERPETIC POLYNEUROPATHY|POSTHERPETIC POLYNEUROPATHY
C2882797|T047|I70.392|ICD10CM|OTHER ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, LEFT LEG|OTH ATHSCL UNSP TYPE BYPASS OF THE EXTREMITIES, LEFT LEG
C0017409|T047|B02.21|ICD10CM|POSTHERPETIC GENICULATE GANGLIONITIS|POSTHERPETIC GENICULATE GANGLIONITIS
C2901807|T047|M86.149|ICD10CM|OTHER ACUTE OSTEOMYELITIS, UNSPECIFIED HAND|OTHER ACUTE OSTEOMYELITIS, UNSPECIFIED HAND
C2842118|T191|C50.529|ICD10CM|MALIGNANT NEOPLASM OF LOWER-OUTER QUADRANT OF UNSPECIFIED MALE BREAST|MALIG NEOPLASM OF LOWER-OUTER QUADRANT OF UNSP MALE BREAST
C2873937|T047|E08.628|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH OTHER SKIN COMPLICATIONS|DIABETES DUE TO UNDERLYING CONDITION W OTH SKIN COMP
C2882798|T047|I70.393|ICD10CM|OTHER ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, BILATERAL LEGS|OTH ATHSCL UNSP TYPE BYPASS OF THE EXTRM, BILATERAL LEGS
C2900495|T047|B02.29|ICD10CM|OTHER POSTHERPETIC NERVOUS SYSTEM INVOLVEMENT|OTHER POSTHERPETIC NERVOUS SYSTEM INVOLVEMENT
C2873935|T047|E08.621|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH FOOT ULCER|DIABETES MELLITUS DUE TO UNDERLYING CONDITION W FOOT ULCER
C2873934|T047|E08.620|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH DIABETIC DERMATITIS|DIABETES DUE TO UNDERLYING CONDITION W DIABETIC DERMATITIS
C2873936|T047|E08.622|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH OTHER SKIN ULCER|DIABETES DUE TO UNDERLYING CONDITION W OTH SKIN ULCER
C2882796|T047|I70.391|ICD10CM|OTHER ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, RIGHT LEG|OTH ATHSCL UNSP TYPE BYPASS OF THE EXTREMITIES, RIGHT LEG
C2888729|T047|L97.521|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF LEFT FOOT LIMITED TO BREAKDOWN OF SKIN|NON-PRS CHRONIC ULCER OTH PRT L FOOT LIMITED TO BRKDWN SKIN
C2888731|T047|L97.523|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF LEFT FOOT WITH NECROSIS OF MUSCLE|NON-PRS CHRONIC ULCER OTH PRT LEFT FOOT W NECROSIS OF MUSCLE
C2888730|T047|L97.522|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF LEFT FOOT WITH FAT LAYER EXPOSED|NON-PRS CHRONIC ULCER OTH PRT LEFT FOOT W FAT LAYER EXPOSED
C4509317|T047|L97.525|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF LEFT FOOT WITH MUSCLE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OTH PRT L FOOT WITH MSL INVL W/O EVD OF NECR
C2888732|T047|L97.524|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF LEFT FOOT WITH NECROSIS OF BONE|NON-PRS CHRONIC ULCER OTH PRT LEFT FOOT W NECROSIS OF BONE
C4509318|T047|L97.526|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF LEFT FOOT WITH BONE INVOLVEMENT WITHOUT EVIDENCE OF NECROSIS|NON-PRS CHR ULC OTH PRT L FOOT WITH BNE INVL W/O EVD OF NECR
C2888733|T047|L97.529|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF LEFT FOOT WITH UNSPECIFIED SEVERITY|NON-PRESSURE CHRONIC ULCER OTH PRT LEFT FOOT W UNSP SEVERITY
C4509319|T047|L97.528|ICD10CM|NON-PRESSURE CHRONIC ULCER OF OTHER PART OF LEFT FOOT WITH OTHER SPECIFIED SEVERITY|NON-PRS CHRONIC ULCER OTH PRT LEFT FOOT WITH OTH SEVERITY
C2859174|T037|S73.014A|ICD10CM|POSTERIOR DISLOCATION OF RIGHT HIP, INITIAL ENCOUNTER|POSTERIOR DISLOCATION OF RIGHT HIP, INITIAL ENCOUNTER
C2883098|T047|I82.421|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF RIGHT ILIAC VEIN|ACUTE EMBOLISM AND THROMBOSIS OF RIGHT ILIAC VEIN
C2883100|T047|I82.423|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF ILIAC VEIN, BILATERAL|ACUTE EMBOLISM AND THROMBOSIS OF ILIAC VEIN, BILATERAL
C2883099|T047|I82.422|ICD10CM|ACUTE EMBOLISM AND THROMBOSIS OF LEFT ILIAC VEIN|ACUTE EMBOLISM AND THROMBOSIS OF LEFT ILIAC VEIN
C2874818|T048|F19.231|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH WITHDRAWAL DELIRIUM|OTH PSYCHOACTIVE SUBSTANCE DEPENDENCE W WITHDRAWAL DELIRIUM
C2874817|T048|F19.230|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH WITHDRAWAL, UNCOMPLICATED|OTH PSYCHOACTIVE SUBSTANCE DEPENDENCE W WITHDRAWAL, UNCOMP
C2874819|T048|F19.232|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE DEPENDENCE WITH WITHDRAWAL WITH PERCEPTUAL DISTURBANCE|OTH PSYCHOACTV SUB DEPEND W W/DRAWAL W PERCEPTL DISTURB
C2889256|T047|M05.469|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSP KNEE
C2855877|T037|S68.113S|ICD10CM|COMPLETE TRAUMATIC METACARPOPHALANGEAL AMPUTATION OF LEFT MIDDLE FINGER, SEQUELA|COMPLETE TRAUMATIC MCP AMPUTATION OF L MID FINGER, SEQUELA
C2889254|T047|M05.461|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT KNEE|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889255|T047|M05.462|ICD10CM|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT KNEE|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT KNEE
C2910915|T033|Z48.21|ICD10CM|ENCOUNTER FOR AFTERCARE FOLLOWING HEART TRANSPLANT|ENCOUNTER FOR AFTERCARE FOLLOWING HEART TRANSPLANT
C2833937|T037|S14.125S|ICD10CM|CENTRAL CORD SYNDROME AT C5 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|CENTRAL CORD SYNDROME AT C5, SEQUELA
C2835818|T037|S24.141A|ICD10CM|BROWN-SEQUARD SYNDROME AT T1 LEVEL OF THORACIC SPINAL CORD, INITIAL ENCOUNTER|BROWN-SEQUARD SYNDROME AT T1, INIT
C2886069|T037|T65.3X2A|ICD10CM|TOXIC EFFECT OF NITRODERIVATIVES AND AMINODERIVATIVES OF BENZENE AND ITS HOMOLOGUES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOX EFF OF NITRODRV/AMINODRV OF BENZN/HOMOLOG, SLF-HRM, INIT
C2833935|T037|S14.125A|ICD10CM|CENTRAL CORD SYNDROME AT C5 LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|CENTRAL CORD SYNDROME AT C5, INIT
C2874228|T047|E70.29|ICD10CM|OTHER DISORDERS OF TYROSINE METABOLISM|OTHER DISORDERS OF TYROSINE METABOLISM
C2833936|T037|S14.125D|ICD10CM|CENTRAL CORD SYNDROME AT C5 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|CENTRAL CORD SYNDROME AT C5, SUBS
C2879948|T037|T48.1X2S|ICD10CM|POISONING BY SKELETAL MUSCLE RELAXANTS [NEUROMUSCULAR BLOCKING AGENTS], INTENTIONAL SELF-HARM, SEQUELA|POISONING BY SKELETAL MUSCLE RELAXANTS, SELF-HARM, SEQUELA
C1879362|T047|E70.21|ICD10CM|TYROSINEMIA|HYPERTYROSINEMIA
C0268482|T047|E70.20|ICD10CM|DISORDER OF TYROSINE METABOLISM, UNSPECIFIED|DISORDER OF TYROSINE METABOLISM, UNSPECIFIED
C2886071|T037|T65.3X2S|ICD10CM|TOXIC EFFECT OF NITRODERIVATIVES AND AMINODERIVATIVES OF BENZENE AND ITS HOMOLOGUES, INTENTIONAL SELF-HARM, SEQUELA|TOX EFF OF NITRODRV/AMINODRV OF BENZN/HOMOLOG, SLF-HRM, SQLA
C2889280|T047|M05.542|ICD10CM|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT HAND|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF LEFT HAND
C2845876|T191|C62.11|ICD10CM|MALIGNANT NEOPLASM OF DESCENDED RIGHT TESTIS|MALIGNANT NEOPLASM OF DESCENDED RIGHT TESTIS
C2845875|T191|C62.10|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED DESCENDED TESTIS|MALIGNANT NEOPLASM OF UNSPECIFIED DESCENDED TESTIS
C2845877|T191|C62.12|ICD10CM|MALIGNANT NEOPLASM OF DESCENDED LEFT TESTIS|MALIGNANT NEOPLASM OF DESCENDED LEFT TESTIS
C2842082|T191|C50.022|ICD10CM|MALIGNANT NEOPLASM OF NIPPLE AND AREOLA, LEFT MALE BREAST|MALIGNANT NEOPLASM OF NIPPLE AND AREOLA, LEFT MALE BREAST
C2889311|T047|M05.642|ICD10CM|RHEUMATOID ARTHRITIS OF LEFT HAND WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF LEFT HAND W INVOLV OF ORGANS AND SYSTEMS
C2838114|T037|S32.434A|ICD10CM|NONDISPLACED FRACTURE OF ANTERIOR COLUMN [ILIOPUBIC] OF RIGHT ACETABULUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP FX OF ANTERIOR COLUMN OF RIGHT ACETABULUM, INIT
C2889312|T047|M05.649|ICD10CM|RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS|RHEU ARTHRITIS OF UNSP HAND W INVOLV OF ORGANS AND SYSTEMS
C2856828|T037|S72.043B|ICD10CM|DISPLACED FRACTURE OF BASE OF NECK OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF BASE OF NK OF UNSP FEMR, INIT FOR OPN FX TYPE I/2
C2856829|T037|S72.043C|ICD10CM|DISPLACED FRACTURE OF BASE OF NECK OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF BASE OF NK OF UNSP FEMR, 7THC
C2856827|T037|S72.043A|ICD10CM|DISPLACED FRACTURE OF BASE OF NECK OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF BASE OF NECK OF UNSP FEMUR, INIT FOR CLOS FX
C2832117|T037|S06.315S|ICD10CM|CONTUSION AND LACERATION OF RIGHT CEREBRUM WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL, SEQUELA|CONTUS/LAC R CEREB W LOC >24 HR W RET CONSC LEV, SEQUELA
C3263930|T046|T84.022A|ICD10CM|INSTABILITY OF INTERNAL RIGHT KNEE PROSTHESIS, INITIAL ENCOUNTER|INSTABILITY OF INTERNAL RIGHT KNEE PROSTHESIS, INIT ENCNTR
C2830409|T033|R40.2314|ICD10CM|COMA SCALE, BEST MOTOR RESPONSE, NONE, 24 HOURS OR MORE AFTER HOSPITAL ADMISSION|COMA SCALE, BEST MOTOR RESPONSE, NONE, 24+HRS
C2830408|T033|R40.2313|ICD10CM|COMA SCALE, BEST MOTOR RESPONSE, NONE, AT HOSPITAL ADMISSION|COMA SCALE, BEST MOTOR RESPONSE, NONE, AT HOSPITAL ADMISSION
C2830407|T033|R40.2312|ICD10CM|COMA SCALE, BEST MOTOR RESPONSE, NONE, AT ARRIVAL TO EMERGENCY DEPARTMENT|COMA SCALE, BEST MOTOR RESPONSE, NONE, EMR
C2830406|T033|R40.2311|ICD10CM|COMA SCALE, BEST MOTOR RESPONSE, NONE, IN THE FIELD [EMT OR AMBULANCE]|COMA SCALE, BEST MOTOR RESPONSE, NONE, IN THE FIELD
C2830405|T033|R40.2310|ICD10CM|COMA SCALE, BEST MOTOR RESPONSE, NONE, UNSPECIFIED TIME|COMA SCALE, BEST MOTOR RESPONSE, NONE, UNSPECIFIED TIME
C0276321|T047|B26.85|ICD10CM|MUMPS ARTHRITIS|MUMPS ARTHRITIS
C2890311|T037|T83.29XA|ICD10CM|OTHER MECHANICAL COMPLICATION OF GRAFT OF URINARY ORGAN, INITIAL ENCOUNTER|MECH COMPL OF GRAFT OF URINARY ORGAN, INITIAL ENCOUNTER
C2900990|T046|M84.451A|ICD10CM|PATHOLOGICAL FRACTURE, RIGHT FEMUR, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, RIGHT FEMUR, INIT ENCNTR FOR FRACTURE
C2902057|T046|M87.246|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED FINGER(S)|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED FINGER(S)
C2902055|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, RIGHT FINGER(S)
C2902056|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, LEFT FINGER(S)
C2902053|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, LEFT HAND
C2902054|T046|M87.243|ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED HAND|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, UNSPECIFIED HAND
C2902052|T046||ICD10CM|OSTEONECROSIS DUE TO PREVIOUS TRAUMA, RIGHT HAND
C2837959|T191|C34.82|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF LEFT BRONCHUS AND LUNG|MALIGNANT NEOPLASM OF OVRLP SITES OF LEFT BRONCHUS AND LUNG
C2837958|T191|C34.81|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF RIGHT BRONCHUS AND LUNG|MALIGNANT NEOPLASM OF OVRLP SITES OF RIGHT BRONCHUS AND LUNG
C2530906|T061|D700|ICD10PCS|CONGENITAL AGRANULOCYTOSIS|RADIATION THERAPY @ LYMPHATIC AND HEMATOLOGIC SYSTEM @ BEAM RADIATION @ BONE MARROW
C2833391|T037|S12.301B|ICD10CM|UNSPECIFIED NONDISPLACED FRACTURE OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP NONDISP FX OF FOURTH CERVICAL VERTEBRA, INIT FOR OPN FX
C2833390|T037|S12.301A|ICD10CM|UNSPECIFIED NONDISPLACED FRACTURE OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP NONDISP FX OF FOURTH CERVICAL VERTEBRA, INIT
C4269440|T037|S02.610A|ICD10CM|FRACTURE OF CONDYLAR PROCESS OF MANDIBLE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FX CONDYLAR PROCESS OF MANDIBLE, UNSPECIFIED SIDE, INIT
C2901017|T046|M84.459A|ICD10CM|PATHOLOGICAL FRACTURE, HIP, UNSPECIFIED, INITIAL ENCOUNTER FOR FRACTURE|PATHOLOGICAL FRACTURE, HIP, UNSP, INIT ENCNTR FOR FRACTURE
C2832360|T037|S06.373S|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF CEREBELLUM WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, SEQUELA|CONTUS/LAC/HEM CRBLM W LOC OF 1-5 HRS 59 MIN, SEQUELA
C2832358|T037|S06.373A|ICD10CM|CONTUSION, LACERATION, AND HEMORRHAGE OF CEREBELLUM WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES, INITIAL ENCOUNTER|CONTUS/LAC/HEM CRBLM W LOC OF 1-5 HRS 59 MIN, INIT
C2889453|T046|M06.349|ICD10CM|RHEUMATOID NODULE, UNSPECIFIED HAND|RHEUMATOID NODULE, UNSPECIFIED HAND
C2889451|T046|M06.341|ICD10CM|RHEUMATOID NODULE, RIGHT HAND|RHEUMATOID NODULE, RIGHT HAND
C2889452|T046|M06.342|ICD10CM|RHEUMATOID NODULE, LEFT HAND|RHEUMATOID NODULE, LEFT HAND
C2835842|T037|S24.151D|ICD10CM|OTHER INCOMPLETE LESION AT T1 LEVEL OF THORACIC SPINAL CORD, SUBSEQUENT ENCOUNTER|OTH INCOMPLETE LESION AT T1, SUBS
C0348364|T191|C46.7|DMDICD10|KAPOSI'S SARCOMA OF OTHER SITES|KAPOSI-SARKOM SONSTIGER LOKALISATIONEN
C2833843|T191|C06.89|ICD10CM|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF OTHER PARTS OF MOUTH|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF OTH PRT MOUTH
C0153563|T191||ICD10CM|KAPOSI'S SARCOMA OF GASTROINTESTINAL SITES
C0153565|T191|C46.3|DMDICD10|KAPOSI'S SARCOMA OF LYMPH NODES|KAPOSI-SARKOM DER LYMPHKNOTEN
C0153562|T191|C46.2|DMDICD10|KAPOSI'S SARCOMA OF PALATE|KAPOSI-SARKOM DES GAUMENS
C2842024|T191|C46.1|ICD10CM|KAPOSI'S SARCOMA OF SOFT TISSUE|KAPOSI'S SARCOMA OF MUSCLE
C0153560|T191|C46.0|DMDICD10|KAPOSI'S SARCOMA OF SKIN|KAPOSI-SARKOM DER HAUT
C4268200|T048|F02.81|ICD10CM|DEMENTIA IN OTHER DISEASES CLASSIFIED ELSEWHERE WITH BEHAVIORAL DISTURBANCE|MAJOR NEUROCOGNITIVE DISORDER IN OTHER DISEASES CLASSIFIED ELSEWHERE WITH VIOLENT BEHAVIOR
C4268197|T048|F02.80|ICD10CM|DEMENTIA IN OTHER DISEASES CLASSIFIED ELSEWHERE WITHOUT BEHAVIORAL DISTURBANCE|MAJOR NEUROCOGNITIVE DISORDER IN OTHER DISEASES CLASSIFIED ELSEWHERE
C0036220|T191|C46.9|DMDICD10|KAPOSI'S SARCOMA, UNSPECIFIED|KAPOSI-SARKOM, NICHT NAEHER BEZEICHNET
C2832696|T037|S06.9X6A|ICD10CM|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, INITIAL ENCOUNTER|UNSP INTCRN INJURY W LOC >24 HR W/O RET CONSC W SURV, INIT
C2835248|T037|S22.028B|ICD10CM|OTHER FRACTURE OF SECOND THORACIC VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH FRACTURE OF SECOND THORACIC VERTEBRA, INIT FOR OPN FX
C2835247|T037|S22.028A|ICD10CM|OTHER FRACTURE OF SECOND THORACIC VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF SECOND THORACIC VERTEBRA, INIT FOR CLOS FX
C2861682|T191|D03.72|ICD10CM|MELANOMA IN SITU OF LEFT LOWER LIMB, INCLUDING HIP|MELANOMA IN SITU OF LEFT LOWER LIMB, INCLUDING HIP
C2882898|T047|I70.549|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF UNSPECIFIED SITE|ATHSCL NONAUT BIO BYPASS OF LEFT LEG W ULCER OF UNSP SITE
C2882897|T047|I70.548|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF OTHER PART OF LOWER LEG|ATHSCL NONAUT BIO BYPASS OF LEFT LEG W ULCER OTH PRT LOW LEG
C2882892|T047|I70.543|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF ANKLE|ATHSCL NONAUT BIO BYPASS OF THE LEFT LEG W ULCER OF ANKLE
C2882891|T047|I70.542|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF CALF|ATHSCL NONAUT BIO BYPASS OF THE LEFT LEG W ULCER OF CALF
C2882890|T047|I70.541|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF THIGH|ATHSCL NONAUT BIO BYPASS OF THE LEFT LEG W ULCER OF THIGH
C2861623|T191||ICD10CM|JUVENILE MYELOMONOCYTIC LEUKEMIA, IN REMISSION
C2882896|T047|I70.545|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF OTHER PART OF FOOT|ATHSCL NONAUT BIO BYPASS OF LEFT LEG W ULCER OTH PRT FOOT
C2882894|T047|I70.544|ICD10CM|ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT(S) OF THE LEFT LEG WITH ULCERATION OF HEEL AND MIDFOOT|ATHSCL NONAUT BIO BYPASS OF LEFT LEG W ULC OF HEEL AND MIDFT
C2885013|T037|T60.0X2S|ICD10CM|TOXIC EFFECT OF ORGANOPHOSPHATE AND CARBAMATE INSECTICIDES, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFF OF ORGANOPHOS AND CARBAMATE INSECT, SLF-HRM, SQLA
C4269403|T037|S02.40DS|ICD10CM|MAXILLARY FRACTURE, LEFT SIDE, SEQUELA|MAXILLARY FRACTURE, LEFT SIDE, SEQUELA
C2874265|T047|E72.8|ICD10CM|OTHER SPECIFIED DISORDERS OF AMINO-ACID METABOLISM|DISORDERS OF BETA-AMINO-ACID METABOLISM
C0002514|T047|E72.9|DMDICD10|DISORDER OF AMINO-ACID METABOLISM, UNSPECIFIED|STOERUNG DES AMINOSAEURESTOFFWECHSELS, NICHT NAEHER BEZEICHNET
C2885011|T037|T60.0X2A|ICD10CM|TOXIC EFFECT OF ORGANOPHOSPHATE AND CARBAMATE INSECTICIDES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFF OF ORGANOPHOS AND CARBAMATE INSECT, SLF-HRM, INIT
C2874190|T047|E23.0|ICD10CM|HYPOPITUITARISM|PITUITARY SHORT STATURE
C1399910|T047||ICD10CM|DISORDERS OF LYSINE AND HYDROXYLYSINE METABOLISM
C0011848|T047|E23.2|DMDICD10|DIABETES INSIPIDUS|DIABETES INSIPIDUS
C0869047|T046|E23.3|DMDICD10|HYPOTHALAMIC DYSFUNCTION, NOT ELSEWHERE CLASSIFIED|HYPOTHALAMISCHE DYSFUNKTION, ANDERENORTS NICHT KLASSIFIZIERT
C4269399|T037|S02.40DB|ICD10CM|MAXILLARY FRACTURE, LEFT SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|MAXILLARY FRACTURE, LEFT SIDE, 7THB
C2874262|T047|E72.4|ICD10CM|DISORDERS OF ORNITHINE METABOLISM|ORNITHINEMIA (TYPES I, II)
C0032002|T047|E23.7|DMDICD10|DISORDER OF PITUITARY GLAND, UNSPECIFIED|STOERUNG DER HYPOPHYSE, NICHT NAEHER BEZEICHNET
C2901909|T047|M86.569|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, UNSPECIFIED TIBIA AND FIBULA|OTH CHRONIC HEMATOGENOUS OSTEOMYELIT, UNSP TIBIA AND FIBULA
C0348992|T047|B38.0|DMDICD10|ACUTE PULMONARY COCCIDIOIDOMYCOSIS|AKUTE KOKZIDIOIDOMYKOSE DER LUNGE
C2901907|T047|M86.561|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, RIGHT TIBIA AND FIBULA|OTH CHRONIC HEMATOGENOUS OSTEOMYELIT, RIGHT TIBIA AND FIBULA
C2901908|T047|M86.562|ICD10CM|OTHER CHRONIC HEMATOGENOUS OSTEOMYELITIS, LEFT TIBIA AND FIBULA|OTH CHRONIC HEMATOGENOUS OSTEOMYELIT, LEFT TIBIA AND FIBULA
C2857496|T037|S72.143A|ICD10CM|DISPLACED INTERTROCHANTERIC FRACTURE OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED INTERTROCHANTERIC FRACTURE OF UNSP FEMUR, INIT
C2882495|T047|I69.133|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING RIGHT NON-DOMINANT SIDE|MONOPLG UPR LMB FOL NTRM INTCRBL HEMOR AFF RIGHT NONDOM SIDE
C2882496|T047|I69.134|ICD10CM|MONOPLEGIA OF UPPER LIMB FOLLOWING NONTRAUMATIC INTRACEREBRAL HEMORRHAGE AFFECTING LEFT NON-DOMINANT SIDE|MONOPLG UPR LMB FOL NTRM INTCRBL HEMOR AFF LEFT NONDOM SIDE
C2838486|T037|S32.699A|ICD10CM|OTHER SPECIFIED FRACTURE OF UNSPECIFIED ISCHIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF UNSP ISCHIUM, INIT FOR CLOS FX
C2889526|T047|M08.011|ICD10CM|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, RIGHT SHOULDER|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS, RIGHT SHOULDER
C2833868|T037|S14.106S|ICD10CM|UNSPECIFIED INJURY AT C6 LEVEL OF CERVICAL SPINAL CORD, SEQUELA|UNSP INJURY AT C6 LEVEL OF CERVICAL SPINAL CORD, SEQUELA
C2888336|T047|L89.144|ICD10CM|PRESSURE ULCER OF LEFT LOWER BACK, STAGE 4|PRESSURE ULCER OF LEFT LOWER BACK, STAGE 4
C2833867|T037|S14.106D|ICD10CM|UNSPECIFIED INJURY AT C6 LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|UNSP INJURY AT C6 LEVEL OF CERVICAL SPINAL CORD, SUBS ENCNTR
C2888324|T047||ICD10CM|PRESSURE ULCER OF LEFT LOWER BACK, UNSTAGEABLE
C2888327|T047|L89.141|ICD10CM|PRESSURE ULCER OF LEFT LOWER BACK, STAGE 1|PRESSURE ULCER OF LEFT LOWER BACK, STAGE 1
C2888330|T047|L89.142|ICD10CM|PRESSURE ULCER OF LEFT LOWER BACK, STAGE 2|PRESSURE ULCER OF LEFT LOWER BACK, STAGE 2
C2888333|T047|L89.143|ICD10CM|PRESSURE ULCER OF LEFT LOWER BACK, STAGE 3|PRESSURE ULCER OF LEFT LOWER BACK, STAGE 3
C2884962|T037|T59.812A|ICD10CM|TOXIC EFFECT OF SMOKE, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF SMOKE, INTENTIONAL SELF-HARM, INIT ENCNTR
C2861618|T191||ICD10CM|ACUTE MONOBLASTIC/MONOCYTIC LEUKEMIA, IN RELAPSE
C2888339|T047|L89.149|ICD10CM|PRESSURE ULCER OF LEFT LOWER BACK, UNSPECIFIED STAGE|PRESSURE ULCER OF LEFT LOWER BACK, UNSPECIFIED STAGE
C3831784|T191|C93.0|ICD10CM|ACUTE MONOBLASTIC/MONOCYTIC LEUKEMIA, NOT HAVING ACHIEVED REMISSION|AML M5
C2861617|T191||ICD10CM|ACUTE MONOBLASTIC/MONOCYTIC LEUKEMIA, IN REMISSION
C2902433|T047|M90.531|ICD10CM|OSTEONECROSIS IN DISEASES CLASSIFIED ELSEWHERE, RIGHT FOREARM|OSTEONECROSIS IN DISEASES CLASSD ELSWHR, RIGHT FOREARM
C2882726|T047|I70.244|ICD10CM|ATHEROSCLEROSIS OF NATIVE ARTERIES OF LEFT LEG WITH ULCERATION OF HEEL AND MIDFOOT|ATHSCL NATIVE ART OF LEFT LEG W ULCER OF HEEL AND MIDFOOT
C0029445|T046|M87.9|DMDICD10|OSTEONECROSIS, UNSPECIFIED|KNOCHENNEKROSE, NICHT NAEHER BEZEICHNET
C2889476|T047|M06.832|ICD10CM|OTHER SPECIFIED RHEUMATOID ARTHRITIS, LEFT WRIST|OTHER SPECIFIED RHEUMATOID ARTHRITIS, LEFT WRIST
C0343898|T047|B39.0|DMDICD10|ACUTE PULMONARY HISTOPLASMOSIS CAPSULATI|AKUTE HISTOPLASMOSE DER LUNGE DURCH HISTOPLASMA CAPSULATUM
C2874844|T048|F19.939|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH WITHDRAWAL, UNSPECIFIED|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSP WITH WITHDRAWAL, UNSP
C2874837|T048|F19.921|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH INTOXICATION WITH DELIRIUM|OTH PSYCHOACTIVE SUBSTANCE USE, UNSP W INTOX W DELIRIUM
C2874843|T048|F19.932|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH WITHDRAWAL WITH PERCEPTUAL DISTURBANCE|OTH PSYCHOACTV SUB USE, UNSP W W/DRAWAL W PERCEPTL DISTURB
C2882398|T047|I63.50|ICD10CM|CEREBRAL INFARCTION DUE TO UNSPECIFIED OCCLUSION OR STENOSIS OF UNSPECIFIED CEREBRAL ARTERY|CEREB INFRC DUE TO UNSP OCCLS OR STENOS OF UNSP CEREB ARTERY
C2874842|T048|F19.931|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH WITHDRAWAL DELIRIUM|OTH PSYCHOACTIVE SUBSTANCE USE, UNSP W WITHDRAWAL DELIRIUM
C4268230|T048|F13.94|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED MOOD DISORDER|SEDATIVE, HYPNOTIC, OR ANXIOLYTIC-INDUCED BIPOLAR OR RELATED DISORDER, WITHOUT USE DISORDER
C2874566|T048|F13.96|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED PERSISTING AMNESTIC DISORDER|SEDATV/HYP/ANXIOLYTC USE, UNSP W PERSIST AMNESTIC DISORDER
C4237402|T048|F13.97|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED PERSISTING DEMENTIA|SEDATIVE, HYPNOTIC, OR ANXIOLYTIC-INDUCED MAJOR NEUROCOGNITIVE DISORDER, WITHOUT USE DISORDER
C2874572|T048|F13.99|ICD10CM|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSPECIFIED WITH UNSPECIFIED SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED DISORDER|SEDATIVE, HYPNOTIC OR ANXIOLYTIC USE, UNSP W UNSP DISORDER
C2833412|T037|S12.34XA|ICD10CM|TYPE III TRAUMATIC SPONDYLOLISTHESIS OF FOURTH CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|TYPE III TRAUM SPONDYLOLYSIS OF FOURTH CERVCAL VERT, INIT
C2890559|T037|T84.091A|ICD10CM|OTHER MECHANICAL COMPLICATION OF INTERNAL LEFT HIP PROSTHESIS, INITIAL ENCOUNTER|MECH COMPL OF INTERNAL LEFT HIP PROSTHESIS, INIT ENCNTR
C4269518|T037|S02.642B|ICD10CM|FRACTURE OF RAMUS OF LEFT MANDIBLE, INITIAL ENCOUNTER FOR OPEN FRACTURE|FRACTURE OF RAMUS OF LEFT MANDIBLE, 7THB
C2889610|T047|M08.839|ICD10CM|OTHER JUVENILE ARTHRITIS, UNSPECIFIED WRIST|OTHER JUVENILE ARTHRITIS, UNSPECIFIED WRIST
C4269517|T037|S02.642A|ICD10CM|FRACTURE OF RAMUS OF LEFT MANDIBLE, INITIAL ENCOUNTER FOR CLOSED FRACTURE|FRACTURE OF RAMUS OF LEFT MANDIBLE, INIT
C2349403|T047||ICD10CM|ACUTE ON CHRONIC GRAFT-VERSUS-HOST DISEASE
C0018133|T047|D89.813|ICD10CM|GRAFT-VERSUS-HOST DISEASE, UNSPECIFIED|GRAFT-VERSUS-HOST DISEASE, UNSPECIFIED
C0856825|T047|D89.810|ICD10CM|ACUTE GRAFT-VERSUS-HOST DISEASE|ACUTE GRAFT-VERSUS-HOST DISEASE
C0867389|T047|D89.811|ICD10CM|CHRONIC GRAFT-VERSUS-HOST DISEASE|CHRONIC GRAFT-VERSUS-HOST DISEASE
C2889608|T047|M08.831|ICD10CM|OTHER JUVENILE ARTHRITIS, RIGHT WRIST|OTHER JUVENILE ARTHRITIS, RIGHT WRIST
C2889609|T047|M08.832|ICD10CM|OTHER JUVENILE ARTHRITIS, LEFT WRIST|OTHER JUVENILE ARTHRITIS, LEFT WRIST
C4269522|T037|S02.642S|ICD10CM|FRACTURE OF RAMUS OF LEFT MANDIBLE, SEQUELA|FRACTURE OF RAMUS OF LEFT MANDIBLE, SEQUELA
C2876185|T037|T32.21|ICD10CM|CORROSIONS INVOLVING 20-29% OF BODY SURFACE WITH 10-19% THIRD DEGREE CORROSION|CORROS 20-29% OF BODY SURFACE W 10-19% THIRD DEGREE CORROS
C2876186|T037|T32.22|ICD10CM|CORROSIONS INVOLVING 20-29% OF BODY SURFACE WITH 20-29% THIRD DEGREE CORROSION|CORROS 20-29% OF BODY SURFACE W 20-29% THIRD DEGREE CORROS
C2883257|T037|T48.992S|ICD10CM|POISONING BY OTHER AGENTS PRIMARILY ACTING ON THE RESPIRATORY SYSTEM, INTENTIONAL SELF-HARM, SEQUELA|POISN BY OTH AGENTS PRIM ACT ON THE RESP SYS, SLF-HRM, SQLA
C4269371|T037|S02.402B|ICD10CM|ZYGOMATIC FRACTURE, UNSPECIFIED SIDE, INITIAL ENCOUNTER FOR OPEN FRACTURE|ZYGOMATIC FRACTURE, UNSPECIFIED SIDE, 7THB
C0338596|T047||ICD10CM|SPASTIC DIPLEGIC CEREBRAL PALSY
C2875323|T019|G80.0|ICD10CM|SPASTIC QUADRIPLEGIC CEREBRAL PALSY|CONGENITAL SPASTIC PARALYSIS (CEREBRAL)
C2889383|T047|M05.879|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED ANKLE AND FOOT|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF UNSP ANK/FT
C0837177|T047|G80.2|ICD10CM|SPASTIC HEMIPLEGIC CEREBRAL PALSY|SPASTIC HEMIPLEGIC CEREBRAL PALSY
C0394005|T047|G80.4|DMDICD10|ATAXIC CEREBRAL PALSY|ATAKTISCHE ZEREBRALPARESE
C0392549|T047|G80.9|DMDICD10|CEREBRAL PALSY, UNSPECIFIED|INFANTILE ZEREBRALPARESE, NICHT NAEHER BEZEICHNET
C2889382|T047|M05.872|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT ANKLE AND FOOT|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF LEFT ANK/FT
C2889381|T047|M05.871|ICD10CM|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT ANKLE AND FOOT|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF RIGHT ANK/FT
C2865547|T037|S88.112D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, LEFT LOWER LEG, SUBSEQUENT ENCOUNTER|COMPLETE TRAUM AMP AT LEV BETW KN AND ANKL, L LOW LEG, SUBS
C2865546|T037|S88.112A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, LEFT LOWER LEG, INITIAL ENCOUNTER|COMPLETE TRAUM AMP AT LEV BETW KN AND ANKL, L LOW LEG, INIT
C2835434|T037|S22.079A|ICD10CM|UNSPECIFIED FRACTURE OF T9-T10 VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF T9-T10 VERTEBRA, INIT FOR CLOS FX
C2835435|T037|S22.079B|ICD10CM|UNSPECIFIED FRACTURE OF T9-T10 VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP FRACTURE OF T9-T10 VERTEBRA, INIT FOR OPN FX
C2832641|T037|S06.892S|ICD10CM|OTHER SPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, SEQUELA|INTCRAN INJ W LOSS OF CONSCIOUSNESS OF 31-59 MIN, SEQUELA
C2865548|T037|S88.112S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION AT LEVEL BETWEEN KNEE AND ANKLE, LEFT LOWER LEG, SEQUELA|COMPLETE TRAUM AMP AT LEV BETW KN AND ANKL, L LOW LEG, SQLA
C2858993|T037|S72.492A|ICD10CM|OTHER FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF LOWER END OF LEFT FEMUR, INIT FOR CLOS FX
C2858994|T037|S72.492B|ICD10CM|OTHER FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|OTH FX LOWER END OF LEFT FEMUR, INIT FOR OPN FX TYPE I/2
C2858995|T037|S72.492C|ICD10CM|OTHER FRACTURE OF LOWER END OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|OTH FX LOWER END OF LEFT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2832639|T037|S06.892A|ICD10CM|OTHER SPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES, INITIAL ENCOUNTER|INTCRAN INJ W LOSS OF CONSCIOUSNESS OF 31-59 MIN, INIT
C4509469|T037|T14.91XS|ICD10CM|SUICIDE ATTEMPT, SEQUELA|SUICIDE ATTEMPT, SEQUELA
C3264402|T047|J84.89|ICD10CM|OTHER SPECIFIED INTERSTITIAL PULMONARY DISEASES|NON-SPECIFIC INTERSTITIAL PNEUMONITIS NOS
C3161107|T047||ICD10CM|SURFACTANT MUTATIONS OF THE LUNG
C3161104|T047|J84.82|ICD10CM|ADULT PULMONARY LANGERHANS CELL HISTIOCYTOSIS|ADULT PLCH
C0751674|T191|J84.81|ICD10CM|LYMPHANGIOLEIOMYOMATOSIS|LYMPHANGIOLEIOMYOMATOSIS
C2878433|T037|T43.292S|ICD10CM|POISONING BY OTHER ANTIDEPRESSANTS, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY OTH ANTIDEPRESSANTS, SELF-HARM, SEQUELA
C2833990|T037|S14.139S|ICD10CM|ANTERIOR CORD SYNDROME AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, SEQUELA|ANT CORD SYNDROME AT UNSP LEVEL OF CERV SPINAL CORD, SEQUELA
C2878046|T037|T42.0X2A|ICD10CM|POISONING BY HYDANTOIN DERIVATIVES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY HYDANTOIN DERIVATIVES, SELF-HARM, INIT
C2857360|T037|S72.131A|ICD10CM|DISPLACED APOPHYSEAL FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED APOPHYSEAL FRACTURE OF RIGHT FEMUR, INIT
C2857361|T037|S72.131B|ICD10CM|DISPLACED APOPHYSEAL FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPLACED APOPHYSEAL FX R FEMUR, INIT FOR OPN FX TYPE I/2
C2857362|T037|S72.131C|ICD10CM|DISPLACED APOPHYSEAL FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPLACED APOPHYSEAL FX R FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2878431|T037|T43.292A|ICD10CM|POISONING BY OTHER ANTIDEPRESSANTS, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY OTH ANTIDEPRESSANTS, SELF-HARM, INIT
C2833988|T037|S14.139A|ICD10CM|ANTERIOR CORD SYNDROME AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, INITIAL ENCOUNTER|ANT CORD SYNDROME AT UNSP LEVEL OF CERV SPINAL CORD, INIT
C2833989|T037|S14.139D|ICD10CM|ANTERIOR CORD SYNDROME AT UNSPECIFIED LEVEL OF CERVICAL SPINAL CORD, SUBSEQUENT ENCOUNTER|ANT CORD SYNDROME AT UNSP LEVEL OF CERV SPINAL CORD, SUBS
C2859115|T037|S72.92XC|ICD10CM|UNSPECIFIED FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|UNSP FRACTURE OF LEFT FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2859113|T037|S72.92XA|ICD10CM|UNSPECIFIED FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF LEFT FEMUR, INIT ENCNTR FOR CLOSED FRACTURE
C2878048|T037|T42.0X2S|ICD10CM|POISONING BY HYDANTOIN DERIVATIVES, INTENTIONAL SELF-HARM, SEQUELA|POISONING BY HYDANTOIN DERIVATIVES, SELF-HARM, SEQUELA
C2857379|T037|S72.132C|ICD10CM|DISPLACED APOPHYSEAL FRACTURE OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPLACED APOPHYSEAL FX L FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2890934|T037|T85.02XA|ICD10CM|DISPLACEMENT OF VENTRICULAR INTRACRANIAL (COMMUNICATING) SHUNT, INITIAL ENCOUNTER|DISPLACEMENT OF VENTRICULAR INTRACRANIAL SHUNT, INIT
C2882746|T047|I70.301|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, RIGHT LEG|UNSP ATHSCL UNSP TYPE BYPASS OF THE EXTREMITIES, RIGHT LEG
C2888929|T047|M01.X11|ICD10CM|DIRECT INFECTION OF RIGHT SHOULDER IN INFECTIOUS AND PARASITIC DISEASES CLASSIFIED ELSEWHERE|DIRECT INFCT OF R SHLDR IN INFEC/PARASTC DIS CLASSD ELSWHR
C2882748|T047|I70.303|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, BILATERAL LEGS|UNSP ATHSCL UNSP TYPE BYPASS OF THE EXTRM, BILATERAL LEGS
C4268403|T047|H40.1124|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, LEFT EYE, INDETERMINATE STAGE|PRIMARY OPEN-ANGLE GLAUCOMA, LEFT EYE, INDETERMINATE STAGE
C4268402|T047|H40.1123|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, LEFT EYE, SEVERE STAGE|PRIMARY OPEN-ANGLE GLAUCOMA, LEFT EYE, SEVERE STAGE
C4268401|T047|H40.1122|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, LEFT EYE, MODERATE STAGE|PRIMARY OPEN-ANGLE GLAUCOMA, LEFT EYE, MODERATE STAGE
C2889185|T047|M05.259|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSP HIP
C4268400|T047|H40.1120|ICD10CM|PRIMARY OPEN-ANGLE GLAUCOMA, LEFT EYE, STAGE UNSPECIFIED|PRIMARY OPEN-ANGLE GLAUCOMA, LEFT EYE, STAGE UNSPECIFIED
C2882750|T047|I70.309|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, UNSPECIFIED EXTREMITY|UNSP ATHSCL UNSP TYPE BYPASS OF THE EXTRM, UNSP EXTREMITY
C2882749|T047|I70.308|ICD10CM|UNSPECIFIED ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT(S) OF THE EXTREMITIES, OTHER EXTREMITY|UNSP ATHSCL UNSP TYPE BYPASS OF THE EXTRM, OTH EXTREMITY
C2889184|T047|M05.252|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT HIP|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT HIP
C2889183|T047|M05.251|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT HIP|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT HIP
C2890525|T037|T84.059A|ICD10CM|PERIPROSTHETIC OSTEOLYSIS OF UNSPECIFIED INTERNAL PROSTHETIC JOINT, INITIAL ENCOUNTER|PERIPROSTH OSTEOLYS OF UNSP INTERNAL PROSTHETIC JOINT, INIT
C2874839|T048|F19.929|ICD10CM|OTHER PSYCHOACTIVE SUBSTANCE USE, UNSPECIFIED WITH INTOXICATION, UNSPECIFIED|OTH PSYCHOACTIVE SUBSTANCE USE, UNSP WITH INTOXICATION, UNSP
C2885305|T037|T63.002A|ICD10CM|TOXIC EFFECT OF UNSPECIFIED SNAKE VENOM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF UNSP SNAKE VENOM, SELF-HARM, INIT
C1719301|T047|B59|ICD10CM|PNEUMOCYSTOSIS|PNEUMONIA DUE TO PNEUMOCYSTIS JIROVECI
C2910363|T019|Q92.61|ICD10CM|MARKER CHROMOSOMES IN NORMAL INDIVIDUAL|MARKER CHROMOSOMES IN NORMAL INDIVIDUAL
C2857789|T037|S72.325C|ICD10CM|NONDISPLACED TRANSVERSE FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|NONDISP TRANSVERSE FX SHAFT OF L FEMR, 7THC
C2889122|T047|M05.051|ICD10CM|FELTY'S SYNDROME, RIGHT HIP|FELTY'S SYNDROME, RIGHT HIP
C2857787|T037|S72.325A|ICD10CM|NONDISPLACED TRANSVERSE FRACTURE OF SHAFT OF LEFT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|NONDISP TRANSVERSE FRACTURE OF SHAFT OF LEFT FEMUR, INIT
C2885307|T037|T63.002S|ICD10CM|TOXIC EFFECT OF UNSPECIFIED SNAKE VENOM, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF UNSP SNAKE VENOM, SELF-HARM, SEQUELA
C2884068|T037|T51.92XA|ICD10CM|TOXIC EFFECT OF UNSPECIFIED ALCOHOL, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF UNSP ALCOHOL, INTENTIONAL SELF-HARM, INIT
C2887778|T047|K50.819|ICD10CM|CROHN'S DISEASE OF BOTH SMALL AND LARGE INTESTINE WITH UNSPECIFIED COMPLICATIONS|CROHN'S DISEASE OF BOTH SMALL AND LG INT W UNSP COMP
C2887777|T047|K50.818|ICD10CM|CROHN'S DISEASE OF BOTH SMALL AND LARGE INTESTINE WITH OTHER COMPLICATION|CROHN'S DISEASE OF BOTH SMALL AND LG INT W OTH COMPLICATION
C2884070|T037|T51.92XS|ICD10CM|TOXIC EFFECT OF UNSPECIFIED ALCOHOL, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF UNSP ALCOHOL, INTENTIONAL SELF-HARM, SEQUELA
C4270189|T046|T83.012A|ICD10CM|BREAKDOWN (MECHANICAL) OF NEPHROSTOMY CATHETER, INITIAL ENCOUNTER|BREAKDOWN (MECHANICAL) OF NEPHROSTOMY CATHETER, INIT
C2887773|T047|K50.811|ICD10CM|CROHN'S DISEASE OF BOTH SMALL AND LARGE INTESTINE WITH RECTAL BLEEDING|CROHN'S DISEASE OF BOTH SMALL AND LG INT W RECTAL BLEEDING
C2887775|T047|K50.813|ICD10CM|CROHN'S DISEASE OF BOTH SMALL AND LARGE INTESTINE WITH FISTULA|CROHN'S DISEASE OF BOTH SMALL AND LARGE INTESTINE W FISTULA
C2887774|T047|K50.812|ICD10CM|CROHN'S DISEASE OF BOTH SMALL AND LARGE INTESTINE WITH INTESTINAL OBSTRUCTION|CROHN'S DISEASE OF BOTH SMALL AND LG INT W INTESTINAL OBST
C2887776|T047|K50.814|ICD10CM|CROHN'S DISEASE OF BOTH SMALL AND LARGE INTESTINE WITH ABSCESS|CROHN'S DISEASE OF BOTH SMALL AND LARGE INTESTINE W ABSCESS
C0349054|T191|C67.8|DMDICD10|MALIGNANT NEOPLASM OF OVERLAPPING SITES OF BLADDER|BOESARTIGE NEUBILDUNG: HARNBLASE, MEHRERE TEILBEREICHE UEBERLAPPEND
C0005684|T191|C67.9|DMDICD10|MALIGNANT NEOPLASM OF BLADDER, UNSPECIFIED|BOESARTIGE NEUBILDUNG: HARNBLASE, NICHT NAEHER BEZEICHNET
C2885269|T037|T62.8X2A|ICD10CM|TOXIC EFFECT OF OTHER SPECIFIED NOXIOUS SUBSTANCES EATEN AS FOOD, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF NOXIOUS SUBSTNC EATEN AS FOOD, SLF-HRM, INIT
C0496828|T191|C67.2|DMDICD10|MALIGNANT NEOPLASM OF LATERAL WALL OF BLADDER|BOESARTIGE NEUBILDUNG: LATERALE HARNBLASENWAND
C0153611|T191|C67.3|DMDICD10|MALIGNANT NEOPLASM OF ANTERIOR WALL OF BLADDER|BOESARTIGE NEUBILDUNG: VORDERE HARNBLASENWAND
C0496826|T191|C67.0|DMDICD10|MALIGNANT NEOPLASM OF TRIGONE OF BLADDER|BOESARTIGE NEUBILDUNG: TRIGONUM VESICAE
C0496827|T191|C67.1|DMDICD10|MALIGNANT NEOPLASM OF DOME OF BLADDER|BOESARTIGE NEUBILDUNG: APEX VESICAE
C0153614|T191|C67.6|DMDICD10|MALIGNANT NEOPLASM OF URETERIC ORIFICE|BOESARTIGE NEUBILDUNG: OSTIUM URETERIS
C0153615|T191|C67.7|DMDICD10|MALIGNANT NEOPLASM OF URACHUS|BOESARTIGE NEUBILDUNG: URACHUS
C0153612|T191|C67.4|DMDICD10|MALIGNANT NEOPLASM OF POSTERIOR WALL OF BLADDER|BOESARTIGE NEUBILDUNG: HINTERE HARNBLASENWAND
C0864965|T191|C67.5|ICD10CM|MALIGNANT NEOPLASM OF BLADDER NECK|MALIGNANT NEOPLASM OF INTERNAL URETHRAL ORIFICE
C2901952|T046|M87.039|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED CARPUS|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED CARPUS
C2901951|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF LEFT CARPUS
C2885271|T037|T62.8X2S|ICD10CM|TOXIC EFFECT OF OTHER SPECIFIED NOXIOUS SUBSTANCES EATEN AS FOOD, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF NOXIOUS SUBSTNC EATEN AS FOOD, SLF-HRM, SQLA
C2901948|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF LEFT ULNA
C2901947|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF RIGHT ULNA
C2901950|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF RIGHT CARPUS
C2901949|T046|M87.036|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED ULNA|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED ULNA
C2901944|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF RIGHT RADIUS
C2901946|T046|M87.033|ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED RADIUS|IDIOPATHIC ASEPTIC NECROSIS OF UNSPECIFIED RADIUS
C2901945|T046||ICD10CM|IDIOPATHIC ASEPTIC NECROSIS OF LEFT RADIUS
C2856049|T037|S68.621S|ICD10CM|PARTIAL TRAUMATIC TRANSPHALANGEAL AMPUTATION OF LEFT INDEX FINGER, SEQUELA|PARTIAL TRAUMATIC TRNSPHAL AMPUTATION OF L IDX FNGR, SEQUELA
C2712816|T056|E002|ICD9CM|CONGENITAL IODINE-DEFICIENCY SYNDROME, MIXED TYPE|ACTIVITIES INVOLVING WATER AND WATER CRAFT
C2712807|T056|E001|ICD9CM|CONGENITAL IODINE-DEFICIENCY SYNDROME, MYXEDEMATOUS TYPE|ACTIVITIES INVOLVING WALKING AND RUNNING
C2712898|T033|E000|ICD9CM|CONGENITAL IODINE-DEFICIENCY SYNDROME, NEUROLOGICAL TYPE|EXTERNAL CAUSE STATUS
C0878801|T033||ICD10CM|ENCOUNTER FOR ADEQUACY TESTING FOR PERITONEAL DIALYSIS
C0878731|T033|Z49.31|ICD10CM|ENCOUNTER FOR ADEQUACY TESTING FOR HEMODIALYSIS|ENCOUNTER FOR ADEQUACY TESTING FOR HEMODIALYSIS
C3165526|T047|E00|DMDICD10|CONGENITAL IODINE-DEFICIENCY SYNDROME, UNSPECIFIED|ANGEBORENES JODMANGELSYNDROM
C2882670|T047|I69.951|ICD10CM|HEMIPLEGIA AND HEMIPARESIS FOLLOWING UNSPECIFIED CEREBROVASCULAR DISEASE AFFECTING RIGHT DOMINANT SIDE|HEMIPLGA FOL UNSP CEREBVASC DISEASE AFF RIGHT DOMINANT SIDE
C2837750|T037|S32.139A|ICD10CM|UNSPECIFIED ZONE III FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP ZONE III FRACTURE OF SACRUM, INIT FOR CLOS FX
C2885077|T037|T60.4X2S|ICD10CM|TOXIC EFFECT OF RODENTICIDES, INTENTIONAL SELF-HARM, SEQUELA|TOXIC EFFECT OF RODENTICIDES, INTENTIONAL SELF-HARM, SEQUELA
C2837751|T037|S32.139B|ICD10CM|UNSPECIFIED ZONE III FRACTURE OF SACRUM, INITIAL ENCOUNTER FOR OPEN FRACTURE|UNSP ZONE III FRACTURE OF SACRUM, INIT FOR OPN FX
C2837882|T037|S32.399A|ICD10CM|OTHER FRACTURE OF UNSPECIFIED ILIUM, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH FRACTURE OF UNSP ILIUM, INIT ENCNTR FOR CLOSED FRACTURE
C2875352|T047|G83.30|ICD10CM|MONOPLEGIA, UNSPECIFIED AFFECTING UNSPECIFIED SIDE|MONOPLEGIA, UNSPECIFIED AFFECTING UNSPECIFIED SIDE
C2875353|T047|G83.31|ICD10CM|MONOPLEGIA, UNSPECIFIED AFFECTING RIGHT DOMINANT SIDE|MONOPLEGIA, UNSPECIFIED AFFECTING RIGHT DOMINANT SIDE
C2875354|T047|G83.32|ICD10CM|MONOPLEGIA, UNSPECIFIED AFFECTING LEFT DOMINANT SIDE|MONOPLEGIA, UNSPECIFIED AFFECTING LEFT DOMINANT SIDE
C2875355|T047|G83.33|ICD10CM|MONOPLEGIA, UNSPECIFIED AFFECTING RIGHT NONDOMINANT SIDE|MONOPLEGIA, UNSPECIFIED AFFECTING RIGHT NONDOMINANT SIDE
C2875356|T047|G83.34|ICD10CM|MONOPLEGIA, UNSPECIFIED AFFECTING LEFT NONDOMINANT SIDE|MONOPLEGIA, UNSPECIFIED AFFECTING LEFT NONDOMINANT SIDE
C0153690|T191|C79.51|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF BONE|SECONDARY MALIGNANT NEOPLASM OF BONE
C0346979|T191|C79.52|ICD10CM|SECONDARY MALIGNANT NEOPLASM OF BONE MARROW|SECONDARY MALIGNANT NEOPLASM OF BONE MARROW
C2889171|T047|M05.222|ICD10CM|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT ELBOW|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2877200|T037|T38.802A|ICD10CM|POISONING BY UNSPECIFIED HORMONES AND SYNTHETIC SUBSTITUTES, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY UNSP HORMONES AND SYNTHETIC SUB, SELF-HARM, INIT
C4268774|T046|M84.754A|ICD10CM|COMPLETE TRANSVERSE ATYPICAL FEMORAL FRACTURE, RIGHT LEG, INITIAL ENCOUNTER FOR FRACTURE|COMPLETE TRANSVERSE ATYP FEMORAL FRACTURE, RIGHT LEG, INIT
C0477404|T047|G71.8|DMDICD10|OTHER PRIMARY DISORDERS OF MUSCLES|SONSTIGE PRIMAERE MYOPATHIEN
C0152936|T047|A20.7|DMDICD10|SEPTICEMIC PLAGUE|PESTSEPSIS
C0524688|T047|A20.2|DMDICD10|PNEUMONIC PLAGUE|LUNGENPEST
C2875337|T184|G81.94|ICD10CM|HEMIPLEGIA, UNSPECIFIED AFFECTING LEFT NONDOMINANT SIDE|HEMIPLEGIA, UNSPECIFIED AFFECTING LEFT NONDOMINANT SIDE
C0375218|T184|G81.90|ICD10CM|HEMIPLEGIA, UNSPECIFIED AFFECTING UNSPECIFIED SIDE|HEMIPLEGIA, UNSPECIFIED AFFECTING UNSPECIFIED SIDE
C2875334|T184|G81.91|ICD10CM|HEMIPLEGIA, UNSPECIFIED AFFECTING RIGHT DOMINANT SIDE|HEMIPLEGIA, UNSPECIFIED AFFECTING RIGHT DOMINANT SIDE
C2875335|T184|G81.92|ICD10CM|HEMIPLEGIA, UNSPECIFIED AFFECTING LEFT DOMINANT SIDE|HEMIPLEGIA, UNSPECIFIED AFFECTING LEFT DOMINANT SIDE
C2875336|T184|G81.93|ICD10CM|HEMIPLEGIA, UNSPECIFIED AFFECTING RIGHT NONDOMINANT SIDE|HEMIPLEGIA, UNSPECIFIED AFFECTING RIGHT NONDOMINANT SIDE
C2910846|T033|Z44.121|ICD10CM|ENCOUNTER FOR FITTING AND ADJUSTMENT OF PARTIAL ARTIFICIAL RIGHT LEG|ENCOUNTER FOR FIT/ADJST OF PARTIAL ARTIFICIAL RIGHT LEG
C2900562|T046|M80.879A|ICD10CM|OTHER OSTEOPOROSIS WITH CURRENT PATHOLOGICAL FRACTURE, UNSPECIFIED ANKLE AND FOOT, INITIAL ENCOUNTER FOR FRACTURE|OTH OSTEOPOR W CURRENT PATH FRACTURE, UNSP ANK/FT, INIT
C4267902|T047|E08.3292|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, LEFT EYE|DIAB WITH MILD NONP RTNOP WITHOUT MACULAR EDEMA, LEFT EYE
C4267903|T047|E08.3293|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, BILATERAL|DIABETES WITH MILD NONP RTNOP WITHOUT MACULAR EDEMA, BI
C4267901|T047|E08.3291|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, RIGHT EYE|DIABETES WITH MILD NONP RTNOP WITHOUT MACULAR EDEMA, R EYE
C4267904|T047|E08.3299|ICD10CM|DIABETES MELLITUS DUE TO UNDERLYING CONDITION WITH MILD NONPROLIFERATIVE DIABETIC RETINOPATHY WITHOUT MACULAR EDEMA, UNSPECIFIED EYE|DIABETES WITH MILD NONP RTNOP WITHOUT MACULAR EDEMA, UNSP
C2869787|T037|S98.112S|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT GREAT TOE, SEQUELA|COMPLETE TRAUMATIC AMPUTATION OF LEFT GREAT TOE, SEQUELA
C2869785|T037|S98.112A|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT GREAT TOE, INITIAL ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF LEFT GREAT TOE, INIT ENCNTR
C2869786|T037|S98.112D|ICD10CM|COMPLETE TRAUMATIC AMPUTATION OF LEFT GREAT TOE, SUBSEQUENT ENCOUNTER|COMPLETE TRAUMATIC AMPUTATION OF LEFT GREAT TOE, SUBS ENCNTR
C2860111|T037|S79.099A|ICD10CM|OTHER PHYSEAL FRACTURE OF UPPER END OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH PHYSEAL FRACTURE OF UPPER END OF UNSP FEMUR, INIT
C2977848|T037|S32.502A|ICD10CM|UNSPECIFIED FRACTURE OF LEFT PUBIS, INITIAL ENCOUNTER FOR CLOSED FRACTURE|UNSP FRACTURE OF LEFT PUBIS, INIT ENCNTR FOR CLOSED FRACTURE
C2831969|T037|S06.0X9S|ICD10CM|CONCUSSION WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION, SEQUELA|CONCUSSION W LOSS OF CONSCIOUSNESS OF UNSP DURATION, SEQUELA
C2883230|T037|T48.902A|ICD10CM|POISONING BY UNSPECIFIED AGENTS PRIMARILY ACTING ON THE RESPIRATORY SYSTEM, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISN BY UNSP AGENTS PRIM ACT ON THE RESP SYS, SLF-HRM, INIT
C0027831|T191||ICD10CM|NEUROFIBROMATOSIS, TYPE 1
C0162678|T191|Q85.00|ICD10CM|NEUROFIBROMATOSIS, UNSPECIFIED|NEUROFIBROMATOSIS, UNSPECIFIED
C1335929|T191|Q85.03|ICD10CM|SCHWANNOMATOSIS|SCHWANNOMATOSIS
C0027832|T191||ICD10CM|NEUROFIBROMATOSIS, TYPE 2
C2902006|T046|M87.144|ICD10CM|OSTEONECROSIS DUE TO DRUGS, RIGHT FINGER(S)|OSTEONECROSIS DUE TO DRUGS, RIGHT FINGER(S)
C2921012|T047|Q85.09|ICD10CM|OTHER NEUROFIBROMATOSIS|OTHER NEUROFIBROMATOSIS
C2883458|T037|T49.7X2S|ICD10CM|POISONING BY DENTAL DRUGS, TOPICALLY APPLIED, INTENTIONAL SELF-HARM, SEQUELA|POISN BY DENTAL DRUGS, TOPICALLY APPLIED, SELF-HARM, SEQUELA
C2883232|T037|T48.902S|ICD10CM|POISONING BY UNSPECIFIED AGENTS PRIMARILY ACTING ON THE RESPIRATORY SYSTEM, INTENTIONAL SELF-HARM, SEQUELA|POISN BY UNSP AGENTS PRIM ACT ON THE RESP SYS, SLF-HRM, SQLA
C2837482|T037|S32.010B|ICD10CM|WEDGE COMPRESSION FRACTURE OF FIRST LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|WEDGE COMPRSN FX FIRST LUM VERTEBRA, INIT FOR OPN FX
C2869855|T037|S98.229A|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF TWO OR MORE UNSPECIFIED LESSER TOES, INITIAL ENCOUNTER|PARTIAL TRAUMATIC AMP OF TWO OR MORE UNSP LESSER TOES, INIT
C2837481|T037|S32.010A|ICD10CM|WEDGE COMPRESSION FRACTURE OF FIRST LUMBAR VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|WEDGE COMPRESSION FRACTURE OF FIRST LUMBAR VERTEBRA, INIT
C2832698|T037|S06.9X6S|ICD10CM|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING, SEQUELA|UNSP INTCRN INJURY W LOC >24 HR W/O RET CONSC W SURV, SQLA
C0838512|T047|M46.39|ICD10CM|INFECTION OF INTERVERTEBRAL DISC (PYOGENIC), MULTIPLE SITES IN SPINE|INFECTION OF INTVRT DISC (PYOGENIC), MULTIPLE SITES IN SPINE
C0838520|T047|M46.38|ICD10CM|INFECTION OF INTERVERTEBRAL DISC (PYOGENIC), SACRAL AND SACROCOCCYGEAL REGION|INFECTION OF INTVRT DISC (PYOGENIC), SACR/SACROCYGL REGION
C0838519|T047|M46.37|ICD10CM|INFECTION OF INTERVERTEBRAL DISC (PYOGENIC), LUMBOSACRAL REGION|INFECTION OF INTVRT DISC (PYOGENIC), LUMBOSACRAL REGION
C0838518|T047|M46.36|ICD10AM|INFECTION OF INTERVERTEBRAL DISC (PYOGENIC), LUMBAR REGION|INFECTION OF INTERVERTEBRAL DISC (PYOGENIC), LUMBAR REGION
C0838517|T047|M46.35|ICD10CM|INFECTION OF INTERVERTEBRAL DISC (PYOGENIC), THORACOLUMBAR REGION|INFECTION OF INTVRT DISC (PYOGENIC), THORACOLUMBAR REGION
C0838516|T047|M46.34|ICD10AM|INFECTION OF INTERVERTEBRAL DISC (PYOGENIC), THORACIC REGION|INFECTION OF INTERVERTEBRAL DISC (PYOGENIC), THORACIC REGION
C0838515|T047|M46.33|ICD10CM|INFECTION OF INTERVERTEBRAL DISC (PYOGENIC), CERVICOTHORACIC REGION|INFECTION OF INTVRT DISC (PYOGENIC), CERVICOTHOR REGION
C0838514|T047|M46.32|ICD10AM|INFECTION OF INTERVERTEBRAL DISC (PYOGENIC), CERVICAL REGION|INFECTION OF INTERVERTEBRAL DISC (PYOGENIC), CERVICAL REGION
C0838513|T047|M46.31|ICD10CM|INFECTION OF INTERVERTEBRAL DISC (PYOGENIC), OCCIPITO-ATLANTO-AXIAL REGION|INFECTION OF INTVRT DISC (PYOGENIC), OCCIPT-ATLAN-AX REGION
C0838512|T047|M46.30|ICD10AM|INFECTION OF INTERVERTEBRAL DISC (PYOGENIC), SITE UNSPECIFIED|INFECTION OF INTERVERTEBRAL DISC (PYOGENIC), MULTIPLE SITES IN SPINE
C2853828|T191|C82.40|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIB, UNSPECIFIED SITE|FOLLICULAR LYMPHOMA GRADE IIIB, UNSPECIFIED SITE
C2853829|T191|C82.41|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIB, LYMPH NODES OF HEAD, FACE, AND NECK|FOLICLAR LYMPHOMA GRADE IIIB, NODES OF HEAD, FACE, AND NECK
C2853830|T191|C82.42|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIB, INTRATHORACIC LYMPH NODES|FOLLICULAR LYMPHOMA GRADE IIIB, INTRATHORACIC LYMPH NODES
C2853831|T191|C82.43|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIB, INTRA-ABDOMINAL LYMPH NODES|FOLLICULAR LYMPHOMA GRADE IIIB, INTRA-ABDOMINAL LYMPH NODES
C2853832|T191|C82.44|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIB, LYMPH NODES OF AXILLA AND UPPER LIMB|FOLICLAR LYMPHOMA GRADE IIIB, NODES OF AXILLA AND UPPER LIMB
C2853833|T191|C82.45|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIB, LYMPH NODES OF INGUINAL REGION AND LOWER LIMB|FOLICLAR LYMPH GRADE IIIB, NODES OF ING RGN AND LOWER LIMB
C2853834|T191|C82.46|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIB, INTRAPELVIC LYMPH NODES|FOLLICULAR LYMPHOMA GRADE IIIB, INTRAPELVIC LYMPH NODES
C2853835|T191|C82.47|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIB, SPLEEN|FOLLICULAR LYMPHOMA GRADE IIIB, SPLEEN
C2853836|T191|C82.48|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIB, LYMPH NODES OF MULTIPLE SITES|FOLLICULAR LYMPHOMA GRADE IIIB, LYMPH NODES MULT SITE
C2853837|T191|C82.49|ICD10CM|FOLLICULAR LYMPHOMA GRADE IIIB, EXTRANODAL AND SOLID ORGAN SITES|FOLICLAR LYMPHOMA GRADE IIIB, EXTRNOD AND SOLID ORGAN SITES
C2854093|T191|C91.12|ICD10CM|CHRONIC LYMPHOCYTIC LEUKEMIA OF B-CELL TYPE IN RELAPSE|CHRONIC LYMPHOCYTIC LEUKEMIA OF B-CELL TYPE IN RELAPSE
C2854092|T191|C91.11|ICD10CM|CHRONIC LYMPHOCYTIC LEUKEMIA OF B-CELL TYPE IN REMISSION|CHRONIC LYMPHOCYTIC LEUKEMIA OF B-CELL TYPE IN REMISSION
C2854091|T191|C91.10|ICD10CM|CHRONIC LYMPHOCYTIC LEUKEMIA OF B-CELL TYPE NOT HAVING ACHIEVED REMISSION|CHRONIC LYMPHOCYTIC LEUK OF B-CELL TYPE NOT ACHIEVE REMIS
C4270513|T046|T85.193A|ICD10CM|OTHER MECHANICAL COMPLICATION OF IMPLANTED ELECTRONIC NEUROSTIMULATOR, GENERATOR, INITIAL ENCOUNTER|MECH COMPL OF IMPLNT ELEC NSTIM, GENERATOR, INIT
C2888830|T047|M00.112|ICD10CM|PNEUMOCOCCAL ARTHRITIS, LEFT SHOULDER|PNEUMOCOCCAL ARTHRITIS, LEFT SHOULDER
C2888829|T047|M00.111|ICD10CM|PNEUMOCOCCAL ARTHRITIS, RIGHT SHOULDER|PNEUMOCOCCAL ARTHRITIS, RIGHT SHOULDER
C2902113|T046|M87.364|ICD10CM|OTHER SECONDARY OSTEONECROSIS, RIGHT FIBULA|OTHER SECONDARY OSTEONECROSIS, RIGHT FIBULA
C2833354|T037|S12.250B|ICD10CM|OTHER TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR OPEN FRACTURE|OTH TRAUM DISPL SPONDYLOLYSIS OF 3RD CERVCAL VERT, 7THB
C2888831|T047|M00.119|ICD10CM|PNEUMOCOCCAL ARTHRITIS, UNSPECIFIED SHOULDER|PNEUMOCOCCAL ARTHRITIS, UNSPECIFIED SHOULDER
C2833353|T037|S12.250A|ICD10CM|OTHER TRAUMATIC DISPLACED SPONDYLOLISTHESIS OF THIRD CERVICAL VERTEBRA, INITIAL ENCOUNTER FOR CLOSED FRACTURE|OTH TRAUM DISPL SPONDYLOLYSIS OF THIRD CERVCAL VERT, INIT
C2869778|T037|S98.029S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION OF UNSPECIFIED FOOT AT ANKLE LEVEL, SEQUELA|PARTIAL TRAUMATIC AMP OF UNSP FOOT AT ANKLE LEVEL, SEQUELA
C4270631|T046|T85.840A|ICD10CM|PAIN DUE TO NERVOUS SYSTEM PROSTHETIC DEVICES, IMPLANTS AND GRAFTS, INITIAL ENCOUNTER|PAIN DUE TO NERVOUS SYSTEM PROSTH DEV/GRFT, INIT
C2854055|T191|C85.91|ICD10CM|NON-HODGKIN LYMPHOMA, UNSPECIFIED, LYMPH NODES OF HEAD, FACE, AND NECK|NON-HODGKIN LYMPHOMA, UNSP, NODES OF HEAD, FACE, AND NECK
C2856620|T037|S72.023A|ICD10CM|DISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISP FX OF EPIPHY (SEPARATION) (UPPER) OF UNSP FEMUR, INIT
C2856621|T037|S72.023B|ICD10CM|DISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISP FX OF EPIPHY (SEPARATION) (UPPER) OF UNSP FEMR, 7THB
C2856622|T037|S72.023C|ICD10CM|DISPLACED FRACTURE OF EPIPHYSIS (SEPARATION) (UPPER) OF UNSPECIFIED FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISP FX OF EPIPHY (SEPARATION) (UPPER) OF UNSP FEMR, 7THC
C2859236|T037|S73.041A|ICD10CM|CENTRAL SUBLUXATION OF RIGHT HIP, INITIAL ENCOUNTER|CENTRAL SUBLUXATION OF RIGHT HIP, INITIAL ENCOUNTER
C2857464|T037|S72.141C|ICD10CM|DISPLACED INTERTROCHANTERIC FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE IIIA, IIIB, OR IIIC|DISPLACED INTERTROCH FX R FEMUR, INIT FOR OPN FX TYPE 3A/B/C
C2857463|T037|S72.141B|ICD10CM|DISPLACED INTERTROCHANTERIC FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR OPEN FRACTURE TYPE I OR II|DISPLACED INTERTROCH FX R FEMUR, INIT FOR OPN FX TYPE I/2
C2857462|T037|S72.141A|ICD10CM|DISPLACED INTERTROCHANTERIC FRACTURE OF RIGHT FEMUR, INITIAL ENCOUNTER FOR CLOSED FRACTURE|DISPLACED INTERTROCHANTERIC FRACTURE OF RIGHT FEMUR, INIT
C2905648|T037|X71.0XXS|ICD10CM|INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION WHILE IN BATHTUB, SEQUELA|INTENTIONAL SELF-HARM BY DROWN WHILE IN BATHTUB, SEQUELA
C2877589|T037|T40.1X2A|ICD10CM|POISONING BY HEROIN, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|POISONING BY HEROIN, INTENTIONAL SELF-HARM, INIT ENCNTR
C2859990|T037|S78.022S|ICD10CM|PARTIAL TRAUMATIC AMPUTATION AT LEFT HIP JOINT, SEQUELA|PARTIAL TRAUMATIC AMPUTATION AT LEFT HIP JOINT, SEQUELA
C2901858|T047|M86.359|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, UNSPECIFIED FEMUR|CHRONIC MULTIFOCAL OSTEOMYELITIS, UNSPECIFIED FEMUR
C2885541|T037|T63.312A|ICD10CM|TOXIC EFFECT OF VENOM OF BLACK WIDOW SPIDER, INTENTIONAL SELF-HARM, INITIAL ENCOUNTER|TOXIC EFFECT OF VENOM OF BLACK WIDOW SPIDER, SELF-HARM, INIT
C2905646|T037|X71.0XXA|ICD10CM|INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION WHILE IN BATHTUB, INITIAL ENCOUNTER|INTENTIONAL SELF-HARM BY DROWN WHILE IN BATHTUB, INIT
C2901857|T047|M86.352|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, LEFT FEMUR|CHRONIC MULTIFOCAL OSTEOMYELITIS, LEFT FEMUR
C2901856|T047|M86.351|ICD10CM|CHRONIC MULTIFOCAL OSTEOMYELITIS, RIGHT FEMUR|CHRONIC MULTIFOCAL OSTEOMYELITIS, RIGHT FEMUR
C2905647|T037|X71.0XXD|ICD10CM|INTENTIONAL SELF-HARM BY DROWNING AND SUBMERSION WHILE IN BATHTUB, SUBSEQUENT ENCOUNTER|INTENTIONAL SELF-HARM BY DROWN WHILE IN BATHTUB, SUBS
C3161109|T047|J84.848|ICD10CM|OTHER INTERSTITIAL  LUNG DISEASES OF CHILDHOOD|OTHER INTERSTITIAL LUNG DISEASES OF CHILDHOOD
C0867812|T037|E896|MTHICD9|POSTPROCEDURAL ADRENOCORTICAL (-MEDULLARY) HYPOFUNCTION|BURNING BY WOOD FIRE IN STOVE OF OTHER BUILDING OR STRUCTURE
C0477305|T047|D55.8|DMDICD10|OTHER ANEMIAS DUE TO ENZYME DISORDERS|SONSTIGE ANAEMIEN DURCH ENZYMDEFEKTE
C0494226|T047|D55|DMDICD10|ANEMIA DUE TO ENZYME DISORDER, UNSPECIFIED|ANAEMIE DURCH ENZYMDEFEKTE
C3161105|T047|J84.841|ICD10CM|NEUROENDOCRINE CELL HYPERPLASIA OF INFANCY|NEUROENDOCRINE CELL HYPERPLASIA OF INFANCY
C3161106|T047|J84.842|ICD10CM|PULMONARY INTERSTITIAL GLYCOGENOSIS|PULMONARY INTERSTITIAL GLYCOGENOSIS
C3161108|T047||ICD10CM|ALVEOLAR CAPILLARY DYSPLASIA WITH VEIN MISALIGNMENT
C2873753|T047|D55.2|ICD10CM|ANEMIA DUE TO DISORDERS OF GLYCOLYTIC ENZYMES|PYRUVATE KINASE [PK] DEFICIENCY ANEMIA
C0475533|T047|D55.3|DMDICD10|ANEMIA DUE TO DISORDERS OF NUCLEOTIDE METABOLISM|ANAEMIE DURCH STOERUNGEN DES NUKLEOTIDSTOFFWECHSELS
C0237987|T047|D55.0|DMDICD10|ANEMIA DUE TO GLUCOSE-6-PHOSPHATE DEHYDROGENASE [G6PD] DEFICIENCY|ANAEMIE DURCH GLUKOSE-6-PHOSPHAT-DEHYDROGENASE[G6PD]-MANGEL
C2873752|T047|D55.1|ICD10CM|ANEMIA DUE TO OTHER DISORDERS OF GLUTATHIONE METABOLISM|ANEMIA (DUE TO) HEMOLYTIC NONSPHEROCYTIC (HEREDITARY), TYPE I
C2845932|T191|C72.30|ICD10CM|MALIGNANT NEOPLASM OF UNSPECIFIED OPTIC NERVE|MALIGNANT NEOPLASM OF UNSPECIFIED OPTIC NERVE
