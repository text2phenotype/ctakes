C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NEUROPATHY|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|CARPAL TUNNEL SYNDROME|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|CARPAL TUNNEL SYNDROMES|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|SYNDROMES, CARPAL TUNNEL|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|SYNDROME, CARPAL TUNNEL|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|CTS (CARPAL TUNNEL SYNDROME)|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|CARPAL TUNNEL SYNDROME |MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|COMPRESSION NEUROPATHY, CARPAL TUNNEL|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|MEDIAN NEUROPATHY, CARPAL TUNNEL|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|CARPAL TUNNEL SYNDROME [DISEASE/FINDING]|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|ENTRAPMENT NEUROPATHY, CARPAL TUNNEL|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|CARPAL TUNNEL SYNDROME, UNSPECIFIED UPPER LIMB|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|AMYOTROPHY, THENAR, OF CARPAL ORIGIN|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|MEDIAN NERVE ENTRAPMENT|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|CARPAL TUNNEL SYNDROME |MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|CTS - CARPAL TUNNEL SYNDROME|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|CTS|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|DISTAL MEDIAN NERVE ENTRAPMENT|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|DISTAL MEDIAN NERVE COMPRESSION|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|MEDIAN NERVE COMPRESSION|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|MEDIAN NERVE ENTRAPMENT |MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|CARPAL TUNNEL; SYNDROME|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|COMPRESSION; MEDIAN NERVE (IN CARPAL TUNNEL)|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|ENTRAPMENT; NEUROPATHIC, NERVE, MEDIAN|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|N.MEDIANUS; COMPRESSION (IN CARPAL TUNNEL)|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|NEUROPATHY; ENTRAPMENT, NERVE, MEDIAN|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|SYNDROME; CARPAL TUNNEL|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|CARPAL TUNNEL MEDIAN NEUROPATHY|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|CARPEL TUNNEL SYNDROME|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0007286|T047|246611002|SNOMEDCT_US|SYNDROME CARPEL TUNNEL|MEDIAN NERVE ENTRAPMENT (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETIC NEUROPATHIES|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|NEUROPATHIES, DIABETIC|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETES WITH NEUROLOGICAL MANIFESTATIONS|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETIC NEUROPATHY|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|NEUROPATHY, DIABETIC|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETIC NEUROPATHIES [DISEASE/FINDING]|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|NEUROPATHY;DIABETIC|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|NEUROPATHY - DIABETIC|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETES + NEUROPATHY|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETIC NEUROPATHY |DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETES MELLITUS WITH NEUROPATHY|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETES MELLITUS WITH NEUROLOGICAL MANIFESTATION|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETES MELLITUS NOS WITH NEUROLOGICAL MANIFESTATION |DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETES MELLITUS NOS WITH NEUROLOGICAL MANIFESTATION|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|NEUROPATHY; DIABETES (MANIFESTATION)|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETIC NEUROPATHY  [AMBIGUOUS]|DIABETIC NEUROPATHY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|FACIAL PARALYSIS|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|PARALYSES, FACIAL|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|PARALYSIS, FACIAL|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|FACIAL PALSIES|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|PALSIES, FACIAL|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|PALSY, FACIAL|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|BELL'S PALSY|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|FACIAL PALSY|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|FACIAL PARALYSIS [DISEASE/FINDING]|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|PALSY;FACIAL|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|FACIAL NERVE PARALYSIS|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|FACIAL NERVE PALSY|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|FACIAL NERVE PALSY (CRANIAL NERVE VII)|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|SEVENTH NERVE PALSY|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|VII NERVE PALSY|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|SEVENTH NERVE PARALYSIS|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|FACIAL NERVE PARALYSIS |FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|FACIAL NERVE PALSIES|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|PARALYSIS OF FACIAL NERVE|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|NERVE PARALYSIS, FACIAL|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|PARALYSIS FACIAL|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|FACIAL PALSY |FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|FACIAL; PARALYSIS|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|PARALYSIS; FACIAL NERVE|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|PARALYSIS; FACIAL|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|FACIAL NERVE PARALYSIS, NOS|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|VII TH NERVE PALSY|FACIAL PALSY (DISORDER)
C0015469|T047|280816001|SNOMEDCT_US|PALSY;VII NERVE|FACIAL PALSY (DISORDER)
C0027813|T047|123254001|SNOMEDCT_US|NEURITIDES|NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|NEURITIS|NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|NEURITIS, NOS|NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|NEURITIS |NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|NEURITIS -RETIRED-|NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|NEURITIDES, PERIPHERAL|NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|PERIPHERAL NEURITIDES|NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|PERIPHERAL NEURITIS|NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|NEURITIS [DISEASE/FINDING]|NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|NEURITIS, PERIPHERAL|NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|NEURITIS;PERIPHERAL|NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|NEURITIS |NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|NEURITIS UNSPECIFIED|NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|NEURITIS UNSPECIFIED |NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|PERIPHERAL NEURITIS NOS|NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|NEURITIS NOS|NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|NEURITIS PERIPHERAL|NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|PERIPHERAL NEURITIS |NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|NEURITIS; PERIPHERAL|NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|PERIPHERAL; NEURITIS|NEURITIS -RETIRED-
C0027813|T047|123254001|SNOMEDCT_US|PERIPHERAL NEURITIS, NOS|NEURITIS -RETIRED-
C0036396|T047|23056005|SNOMEDCT_US|SCIATICA|SCIATICA (DISORDER)
C0036396|T047|23056005|SNOMEDCT_US|SCIATICA |SCIATICA (DISORDER)
C0036396|T047|23056005|SNOMEDCT_US|ISCHIAS|SCIATICA (DISORDER)
C0036396|T047|23056005|SNOMEDCT_US|NEURALGIAS, SCIATIC|SCIATICA (DISORDER)
C0036396|T047|23056005|SNOMEDCT_US|SCIATIC NEURALGIAS|SCIATICA (DISORDER)
C0036396|T047|23056005|SNOMEDCT_US|SCIATICA, UNSPECIFIED SIDE|SCIATICA (DISORDER)
C0036396|T047|23056005|SNOMEDCT_US|SCIATIC NEURALGIA|SCIATICA (DISORDER)
C0036396|T047|23056005|SNOMEDCT_US|SCIATICA [DISEASE/FINDING]|SCIATICA (DISORDER)
C0036396|T047|23056005|SNOMEDCT_US|NEURALGIA, SCIATIC|SCIATICA (DISORDER)
C0036396|T047|23056005|SNOMEDCT_US|SCIATIA|SCIATICA (DISORDER)
C0036396|T047|23056005|SNOMEDCT_US|SCIATICA |SCIATICA (DISORDER)
C0036396|T047|23056005|SNOMEDCT_US|ISCHIALGIA|SCIATICA (DISORDER)
C0036396|T047|23056005|SNOMEDCT_US|COTUGNO'S DISEASE|SCIATICA (DISORDER)
C0036396|T047|23056005|SNOMEDCT_US|NEURALGIA-NEURITIS OF SCIATIC NERVE|SCIATICA (DISORDER)
C0036396|T047|23056005|SNOMEDCT_US|SCIATICA NEURALGIA|SCIATICA (DISORDER)
C0036396|T047|23056005|SNOMEDCT_US|NEURALGIA OR NEURITIS OF SCIATIC NERVE|SCIATICA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|FOTHERGILL'S NEURALGIA|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|NEURALGIAS, TRIGEMINAL|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TRIGEMINAL NEURALGIA|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TRIGEMINAL NEURALGIAS|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|NEURALGIA, TRIGEMINAL|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|FOTHERGILL DIS|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TIC DOULOUREUX|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TRIFOCAL NEURALGIA|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TIC DOLOREUX|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|DISEASE, FOTHERGILL|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|NEURALGIA, EPILEPTIFORM|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|EPILEPTIFORM NEURALGIAS|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|NEURALGIAS, EPILEPTIFORM|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|NEURALGIA, TRIFACIAL|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|NEURALGIAS, TRIFACIAL|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TRIFACIAL NEURALGIAS|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|FOTHERGILL DISEASE|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TRIFACIAL NEURALGIA|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TRIGEMINAL NEURALGIA [DISEASE/FINDING]|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|EPILEPTIFORM NEURALGIA|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TIC DOULEUREUX|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TRIGEMINAL NEURALGIA NOS|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TRIGEMINAL NEURALGIA [NO DRUGS HERE] |TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TRIGEMINAL NEURALGIA [NO DRUGS HERE]|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TRIGEMINAL NEURALGIA NOS |TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TRIGEMINAL NEURALGIA |TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TRIGEMINAL NEURALGIA |TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|NEURALGIA TRIGEMINAL|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TN - TRIGEMINAL NEURALGIA|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|FOTHERGILL; NEURALGIA|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|FOTHERGILL; TRIGEMINAL NEURALGIA|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|DOULOUREUX; TIC|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|NEURALGIA; FOTHERGILL|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|NEURALGIA; CRANIAL NERVE, FIFTH OR TRIGEMINAL|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|NEURALGIA; TRIFACIAL|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|NEURALGIA; TRIGEMINAL|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|PAIN; TRIGEMINAL|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TIC; DOULOUREUX|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TRIFACIAL; NEURALGIA|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TRIGEMINAL NEURALGIA; FOTHERGILL|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TRIGEMINAL; NEURALGIA|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TRIGEMINAL; PAIN|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TRIGEMINAL NEURALGIA, NOS|TRIGEMINAL NEURALGIA (DISORDER)
C0040997|T047|31681005|SNOMEDCT_US|TIC DOLOUREUX|TRIGEMINAL NEURALGIA (DISORDER)
C0596694|T047||SNOMEDCT_US|HEREDITARY PERIPHERAL NERVOUS SYSTEM DISORDER
C0151313|T047|95662005|SNOMEDCT_US|PERIPHERAL SENSORY NEUROPATHY|SENSORY NEUROPATHY (DISORDER)
C0151313|T047|95662005|SNOMEDCT_US|SENSORY NEUROPATHY|SENSORY NEUROPATHY (DISORDER)
C0151313|T047|95662005|SNOMEDCT_US|PERIPHERAL NEUROPATHY, SENSORY|SENSORY NEUROPATHY (DISORDER)
C0151313|T047|95662005|SNOMEDCT_US|SENSORY PERIPHERAL NEUROPATHIES|SENSORY NEUROPATHY (DISORDER)
C0151313|T047|95662005|SNOMEDCT_US|SENSORY PERIPHERAL NEUROPATHY|SENSORY NEUROPATHY (DISORDER)
C0151313|T047|95662005|SNOMEDCT_US|SENSORY NEUROPATHY |SENSORY NEUROPATHY (DISORDER)
C0027796|T047|123253007|SNOMEDCT_US|SLIGHTY MORE SPECIFIC FOR PERIPHERAL NEUROPATHY, SO INCLUDING THESE|NEURALGIA -RETIRED-
C0027796|T047|123253007|SNOMEDCT_US|PAIN, NEUROPATHIC|NEURALGIA -RETIRED-
C0027796|T047|123253007|SNOMEDCT_US|NEUROPATHIC PAIN|NEURALGIA -RETIRED-
C0235025|T047|95663000|SNOMEDCT_US|PERIPHERAL MOTOR NEUROPATHY|PERIPHERAL MOTOR NEUROPATHY (DISORDER)
C0235025|T047|95663000|SNOMEDCT_US|MOTOR NEUROPATHY|PERIPHERAL MOTOR NEUROPATHY (DISORDER)
C0235025|T047|95663000|SNOMEDCT_US|MOTOR NEURITIDES|PERIPHERAL MOTOR NEUROPATHY (DISORDER)
C0235025|T047|95663000|SNOMEDCT_US|MOTOR NEURITIS|PERIPHERAL MOTOR NEUROPATHY (DISORDER)
C0235025|T047|95663000|SNOMEDCT_US|NEURITIDES, MOTOR|PERIPHERAL MOTOR NEUROPATHY (DISORDER)
C0235025|T047|95663000|SNOMEDCT_US|MOTOR PERIPHERAL NEUROPATHY|PERIPHERAL MOTOR NEUROPATHY (DISORDER)
C0235025|T047|95663000|SNOMEDCT_US|NEURITIS MOTOR|PERIPHERAL MOTOR NEUROPATHY (DISORDER)
C0235025|T047|95663000|SNOMEDCT_US|NEURITIS, MOTOR|PERIPHERAL MOTOR NEUROPATHY (DISORDER)
C0235025|T047|95663000|SNOMEDCT_US|PERIPHERAL MOTOR NEUROPATHY |PERIPHERAL MOTOR NEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOLIC POLYNEUROPATHY|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL IND POLYNEUROPATHY|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL IND PERIPHERAL NEUROPATHY|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|PERIPHERAL NEUROPATHY ALCOHOL IND|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL RELAT POLYNEUROPATHY|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL RELAT AUTONOMIC POLYNEUROPATHY|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL-INDUCED POLYNEUROPATHY -RETIRED-|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOLIC POLYNEUROPATHY |ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|POLYNEUROPATHY ALCOHOLIC|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL-RELATED AUTONOMIC POLYNEUROPATHIES|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|AUTONOMIC POLYNEUROPATHIES, ALCOHOL-RELATED|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|POLYNEUROPATHIES, ALCOHOL-RELATED AUTONOMIC|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL RELATED AUTONOMIC POLYNEUROPATHY|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|AUTONOMIC POLYNEUROPATHY, ALCOHOL-RELATED|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|POLYNEUROPATHY, ALCOHOL-RELATED AUTONOMIC|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL INDUCED PERIPHERAL NEUROPATHY|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL-INDUCED PERIPHERAL NEUROPATHIES|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|NEUROPATHIES, ALCOHOL-INDUCED PERIPHERAL|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|NEUROPATHY, ALCOHOL-INDUCED PERIPHERAL|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|PERIPHERAL NEUROPATHIES, ALCOHOL-INDUCED|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|PERIPHERAL NEUROPATHY, ALCOHOL INDUCED|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL-INDUCED POLYNEUROPATHIES|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|POLYNEUROPATHIES, ALCOHOL-INDUCED|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL INDUCED POLYNEUROPATHY|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|POLYNEUROPATHY, ALCOHOL-INDUCED|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL-RELATED POLYNEUROPATHIES|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|POLYNEUROPATHIES, ALCOHOL-RELATED|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL RELATED POLYNEUROPATHY|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|POLYNEUROPATHY, ALCOHOL-RELATED|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOLIC NEUROPATHIES|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOLIC NEUROPATHY|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|NEUROPATHIES, ALCOHOLIC|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOLIC POLYNEURITIDES|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOLIC POLYNEURITIS|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|POLYNEURITIDES, ALCOHOLIC|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOLIC POLYNEUROPATHIES|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|POLYNEUROPATHIES, ALCOHOLIC|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|NEUROPATHY, ALCOHOLIC|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|POLYNEURITIS, ALCOHOLIC|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|POLYNEUROPATHY, ALCOHOLIC|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOLIC NEUROPATHY [DISEASE/FINDING]|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL-INDUCED PERIPHERAL NEUROPATHY|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL-INDUCED POLYNEUROPATHY|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|PERIPHERAL NEUROPATHY, ALCOHOL-INDUCED|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL-RELATED AUTONOMIC POLYNEUROPATHY|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL-RELATED POLYNEUROPATHY|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|NEUROPATHY;ALCOHOLIC|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL-INDUCED POLYNEUROPATHY |ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL-RELATED POLYNEUROPATHY |ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOLIC PERIPHERAL NEUROPATHY|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOLIC POLYNEUROPATHY |ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|POLYNEUROPATHY; ALCOHOLIC|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|POLYNEUROPATHY; ALCOHOL|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0085677|T047|123050003|SNOMEDCT_US|ALCOHOL; POLYNEUROPATHY|ALCOHOL-INDUCED POLYNEUROPATHY (DISORDER)
C0393842|T047||SNOMEDCT_US|POLYNEUROPATHY IN NEOPLASTIC DISEASE
C0393842|T047||SNOMEDCT_US|MALIGNANT NEOPLASM; POLYNEUROPATHY (ETIOLOGY)
C0393842|T047||SNOMEDCT_US|MALIGNANT NEOPLASM; POLYNEUROPATHY (MANIFESTATION)
C0393842|T047||SNOMEDCT_US|NEOPLASM; POLYNEUROPATHY (MANIFESTATION)
C0393842|T047||SNOMEDCT_US|POLYNEUROPATHY; MALIGNANT NEOPLASM (ETIOLOGY)
C0393842|T047||SNOMEDCT_US|POLYNEUROPATHY; MALIGNANT NEOPLASM (MANIFESTATION)
C0393842|T047||SNOMEDCT_US|POLYNEUROPATHY; NEOPLASM (MANIFESTATION)
C0270932|T047|77659000|SNOMEDCT_US|POLYNEUROPATHY IN MALIGNANT DISEASE|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|PERIPHERAL NEUROPATHY PARANEOPL|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|PARANEOPL POLYNEUROPATHY|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|NEUROPATHY PARANEOPL|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|POLYNEUROPATHY PARANEOPL|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|PARANEOPL PERIPHERAL NEUROPATHY|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|PARANEOPL NEUROPATHY|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|POLYNEUROPATHY DUE TO MALIGNANT DISEASE |PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|POLYNEUROPATHY DUE TO MALIGNANT DISEASE|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|NEUROPATHIES, PARANEOPLASTIC|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|PARANEOPLASTIC NEUROPATHIES|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|NEUROPATHIES, PARANEOPLASTIC PERIPHERAL|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|NEUROPATHY, PARANEOPLASTIC PERIPHERAL|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|PARANEOPLASTIC PERIPHERAL NEUROPATHIES|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|PERIPHERAL NEUROPATHIES, PARANEOPLASTIC|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|PARANEOPLASTIC POLYNEUROPATHIES|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|POLYNEUROPATHIES, PARANEOPLASTIC|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|PARANEOPLASTIC POLYNEUROPATHY|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|NEUROPATHY IN MALIG DIS|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|PARANEOPLASTIC NEUROPATHY|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|NEUROPATHY, PARANEOPLASTIC|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|PARANEOPLASTIC PERIPHERAL NEUROPATHY|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|POLYNEUROPATHY, PARANEOPLASTIC|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|PARANEOPLASTIC POLYNEUROPATHY [DISEASE/FINDING]|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|PERIPHERAL NEUROPATHY, PARANEOPLASTIC|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|PARANEOPLASTIC PERIPHERAL NEUROPATHY |PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|CARCINOMATOUS NEUROPATHY|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|POLYNEUROPATHY IN MALIGNANCY|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|CARCINOMATOUS PERIPHERAL NEUROPATHY|PARANEOPLASTIC NEUROPATHY (DISORDER)
C0270932|T047|77659000|SNOMEDCT_US|PARANEOPLASTIC NEUROPATHY |PARANEOPLASTIC NEUROPATHY (DISORDER)
C0859672|T047||SNOMEDCT_US|OTHER HEREDITARY AND IDIOPATHIC PERIPHERAL NEUROPATHY
C0859672|T047||SNOMEDCT_US|HEREDITARY AND IDIOPATHIC PERIPHERAL NEUROPATHY, OTHER
C0859673|T047||SNOMEDCT_US|UNSPECIFIED HEREDITARY AND IDIOPATHIC PERIPHERAL NEUROPATHY
C0859673|T047||SNOMEDCT_US|IDIO PERIPH NEURPTHY NOS
C0477394|T047|194520003|SNOMEDCT_US|OTHER SPECIFIED POLYNEUROPATHIES|[X]OTHER SPECIFIED POLYNEUROPATHIES (DISORDER)
C0477394|T047|194520003|SNOMEDCT_US|[X]OTHER SPECIFIED POLYNEUROPATHIES|[X]OTHER SPECIFIED POLYNEUROPATHIES (DISORDER)
C0477394|T047|194520003|SNOMEDCT_US|[X]OTHER SPECIFIED POLYNEUROPATHIES |[X]OTHER SPECIFIED POLYNEUROPATHIES (DISORDER)
C0494489|T047|609592007|SNOMEDCT_US|MONONEUROPATHIES OF LOWER LIMB|MONONEUROPATHY OF LOWER LIMB (DISORDER)
C0494489|T047|609592007|SNOMEDCT_US|MONONEUROPATHY OF LOWER LIMB, UNSPECIFIED|MONONEUROPATHY OF LOWER LIMB (DISORDER)
C0494489|T047|609592007|SNOMEDCT_US|UNSPECIFIED MONONEUROPATHY OF UNSPECIFIED LOWER LIMB|MONONEUROPATHY OF LOWER LIMB (DISORDER)
C0494489|T047|609592007|SNOMEDCT_US|UNSPECIFIED MONONEUROPATHY OF LOWER LIMB|MONONEUROPATHY OF LOWER LIMB (DISORDER)
C0494489|T047|609592007|SNOMEDCT_US|MONONEUROPATHY OF LOWER LIMB |MONONEUROPATHY OF LOWER LIMB (DISORDER)
C0494489|T047|609592007|SNOMEDCT_US|MONONEUROPATHY OF LOWER LIMB|MONONEUROPATHY OF LOWER LIMB (DISORDER)
C0154762|T047|7339009|SNOMEDCT_US|POLYNEUROPATHY DUE TO DRUGS|POLYNEUROPATHY DUE TO DRUG (DISORDER)
C0154762|T047|7339009|SNOMEDCT_US|DRUG-INDUCED POLYNEUROPATHY|POLYNEUROPATHY DUE TO DRUG (DISORDER)
C0154762|T047|7339009|SNOMEDCT_US|DRUG-INDUCED POLYNEUROPATHY |POLYNEUROPATHY DUE TO DRUG (DISORDER)
C0154762|T047|7339009|SNOMEDCT_US|NEUROPATHY DUE TO DRUGS|POLYNEUROPATHY DUE TO DRUG (DISORDER)
C0154762|T047|7339009|SNOMEDCT_US|POLYNEUROPATHY DUE TO DRUG |POLYNEUROPATHY DUE TO DRUG (DISORDER)
C0154762|T047|7339009|SNOMEDCT_US|POLYNEUROPATHY CAUSED BY DRUG |POLYNEUROPATHY DUE TO DRUG (DISORDER)
C0154762|T047|7339009|SNOMEDCT_US|POLYNEUROPATHY CAUSED BY DRUG|POLYNEUROPATHY DUE TO DRUG (DISORDER)
C0154762|T047|7339009|SNOMEDCT_US|DRUG-RELATED POLYNEUROPATHY|POLYNEUROPATHY DUE TO DRUG (DISORDER)
C0154762|T047|7339009|SNOMEDCT_US|POLYNEUROPATHY DUE TO DRUG|POLYNEUROPATHY DUE TO DRUG (DISORDER)
C0154762|T047|7339009|SNOMEDCT_US|POLYNEUROPATHY DUE TO DRUG, NOS|POLYNEUROPATHY DUE TO DRUG (DISORDER)
C0494518|T047||SNOMEDCT_US|AUTONOMIC NEUROPATHY IN ENDOCRINE AND METABOLIC DISEASES
C0494518|T047||SNOMEDCT_US|NEUROPATHY; PERIPHERAL, AUTONOMIC, IN METABOLIC DISEASE (MANIFESTATION)
C0235023|T047||SNOMEDCT_US|NEURITIS BULBAR
C0235026|T047||SNOMEDCT_US|NEURITIDES, SENSORY
C0235026|T047||SNOMEDCT_US|SENSORY NEURITIDES
C0235026|T047||SNOMEDCT_US|SENSORY NEURITIS
C0235026|T047||SNOMEDCT_US|NEURITIS SENSORY
C0235026|T047||SNOMEDCT_US|NEURITIS, SENSORY
C0235919|T047||SNOMEDCT_US|NERVE ROOT LIAISON
C0235919|T047||SNOMEDCT_US|NERVE ROOT LESION
C0235919|T047||SNOMEDCT_US|NERVE ROOT LESION NOS
C0238309|T047|129611009|SNOMEDCT_US|ISCHAEMIC NEUROPATHY|ISCHEMIC PERIPHERAL NEUROPATHY (DISORDER)
C0238309|T047|129611009|SNOMEDCT_US|ISCHEMIC NEUROPATHY|ISCHEMIC PERIPHERAL NEUROPATHY (DISORDER)
C0238309|T047|129611009|SNOMEDCT_US|ISCHAEMIC PERIPHERAL NEUROPATHY|ISCHEMIC PERIPHERAL NEUROPATHY (DISORDER)
C0238309|T047|129611009|SNOMEDCT_US|ISCHEMIC NEUROPATHY |ISCHEMIC PERIPHERAL NEUROPATHY (DISORDER)
C0238309|T047|129611009|SNOMEDCT_US|ISCHEMIC PERIPHERAL NEUROPATHY |ISCHEMIC PERIPHERAL NEUROPATHY (DISORDER)
C0238309|T047|129611009|SNOMEDCT_US|ISCHEMIC PERIPHERAL NEUROPATHY|ISCHEMIC PERIPHERAL NEUROPATHY (DISORDER)
C0393807|T047|128203003|SNOMEDCT_US|CMT6|HMSN VI
C0393807|T047|128203003|SNOMEDCT_US|HEREDITARY MOTOR AND SENSORY NEUROPATHY WITH OPTIC ATROPHY |HMSN VI
C0393807|T047|128203003|SNOMEDCT_US|HMSN VI|HMSN VI
C0393807|T047|128203003|SNOMEDCT_US|PERIPHERAL NEUROPATHY AND OPTIC ATROPHY|HMSN VI
C0393807|T047|128203003|SNOMEDCT_US|CHARCOT-MARIE-TOOTH DISEASE, TYPE 6|HMSN VI
C0393807|T047|128203003|SNOMEDCT_US|HMSN6|HMSN VI
C0393807|T047|128203003|SNOMEDCT_US|HEREDITARY MOTOR AND SENSORY NEUROPATHY VI|HMSN VI
C0393807|T047|128203003|SNOMEDCT_US|HEREDITARY MOTOR AND SENSORY NEUROPATHY WITH OPTIC ATROPHY|HMSN VI
C0393807|T047|128203003|SNOMEDCT_US|HEREDITARY MOTOR AND SENSORY NEUROPATHY WITH OPTIC ATROPHY |HMSN VI
C0393807|T047|128203003|SNOMEDCT_US|NEUROPATHY, HEREDITARY MOTOR AND SENSORY, TYPE VI|HMSN VI
C0393807|T047|128203003|SNOMEDCT_US|HSMN6|HMSN VI
C0393807|T047|128203003|SNOMEDCT_US|HEREDITARY MOTOR AND SENSORY NEUROPATHY TYPE VI|HMSN VI
C0393807|T047|128203003|SNOMEDCT_US|HEREDITARY MOTOR-SENSORY NEUROPATHY WITH OPTIC ATROPHY|HMSN VI
C0393807|T047|128203003|SNOMEDCT_US|HEREDITARY MOTOR-SENSORY NEUROPATHY, TYPE VI|HMSN VI
C0393807|T047|128203003|SNOMEDCT_US|HEREDITARY SENSORY AND MOTOR NEUROPATHY, TYPE VI|HMSN VI
C0392553|T047|65017003|SNOMEDCT_US|HEREDITARY PERIPHERAL NEUROPATHY |HEREDITARY PERIPHERAL NEUROPATHY (DISORDER)
C0392553|T047|65017003|SNOMEDCT_US|HEREDITARY PERIPHERAL NEUROPATHY|HEREDITARY PERIPHERAL NEUROPATHY (DISORDER)
C0392553|T047|65017003|SNOMEDCT_US|HERED PERIPH NEUROPATHY|HEREDITARY PERIPHERAL NEUROPATHY (DISORDER)
C0392553|T047|65017003|SNOMEDCT_US|HEREDITARY PERIPHERAL NEUROPATHY NOS|HEREDITARY PERIPHERAL NEUROPATHY (DISORDER)
C0392553|T047|65017003|SNOMEDCT_US|HEREDITARY PERIPHERAL NEUROPATHY NOS |HEREDITARY PERIPHERAL NEUROPATHY (DISORDER)
C0392553|T047|65017003|SNOMEDCT_US|PERIPHERAL NEUROPATHY HEREDITARY|HEREDITARY PERIPHERAL NEUROPATHY (DISORDER)
C0392553|T047|65017003|SNOMEDCT_US|HEREDITARY PERIPHERAL NEUROPATHY |HEREDITARY PERIPHERAL NEUROPATHY (DISORDER)
C0392553|T047|65017003|SNOMEDCT_US|HEREDITARY PERIPHERAL NEUROPATHY, NOS|HEREDITARY PERIPHERAL NEUROPATHY (DISORDER)
C0154690|T047|86489003|SNOMEDCT_US|IDIOPATHIC PERIPHERAL AUTONOMIC NEUROPATHY|IDIOPATHIC PERIPHERAL AUTONOMIC NEUROPATHY (DISORDER)
C0154690|T047|86489003|SNOMEDCT_US|IDIOPATHIC PERIPHERAL AUTONOMIC NEUROPATHY |IDIOPATHIC PERIPHERAL AUTONOMIC NEUROPATHY (DISORDER)
C0154690|T047|86489003|SNOMEDCT_US|IDIOPATHIC PERIPHERAL AUTONOMIC NEUROPATHY NOS|IDIOPATHIC PERIPHERAL AUTONOMIC NEUROPATHY (DISORDER)
C0154690|T047|86489003|SNOMEDCT_US|IDIOPATHIC PERIPHERAL AUTONOMIC NEUROPATHY |IDIOPATHIC PERIPHERAL AUTONOMIC NEUROPATHY (DISORDER)
C0154690|T047|86489003|SNOMEDCT_US|IDIOPATHIC PERIPHERAL AUTONOMIC NEUROPATHY NOS |IDIOPATHIC PERIPHERAL AUTONOMIC NEUROPATHY (DISORDER)
C0154690|T047|86489003|SNOMEDCT_US|NEUROPATHY; PERIPHERAL, AUTONOMIC, IDIOPATHIC|IDIOPATHIC PERIPHERAL AUTONOMIC NEUROPATHY (DISORDER)
C0154754|T047|193157005|SNOMEDCT_US|HEREDITARY AND IDIOPATHIC PERIPHERAL NEUROPATHY|HEREDITARY AND IDIOPATHIC PERIPHERAL NEUROPATHY (DISORDER)
C0154754|T047|193157005|SNOMEDCT_US|HEREDITARY AND IDIOPATHIC NEUROPATHY|HEREDITARY AND IDIOPATHIC PERIPHERAL NEUROPATHY (DISORDER)
C0154754|T047|193157005|SNOMEDCT_US|HEREDITARY AND IDIOPATHIC NEUROPATHY, UNSPECIFIED|HEREDITARY AND IDIOPATHIC PERIPHERAL NEUROPATHY (DISORDER)
C0154754|T047|193157005|SNOMEDCT_US|HEREDITARY AND IDIOPATHIC PERIPHERAL NEUROPATHY |HEREDITARY AND IDIOPATHIC PERIPHERAL NEUROPATHY (DISORDER)
C0154691|T047||SNOMEDCT_US|PERIPHERAL AUTONOMIC NEUROPATHY IN DISORDERS CLASSIFIED ELSEWHERE
C0154691|T047||SNOMEDCT_US|AUT NEUROPTHY IN OTH DIS
C0154757|T047||SNOMEDCT_US|OTHER SPECIFIED IDIOPATHIC PERIPHERAL NEUROPATHY
C0154757|T047||SNOMEDCT_US|IDIO PERIPH NEURPTHY NEC
C0041848|T047||SNOMEDCT_US|UNSPECIFIED IDIOPATHIC PERIPHERAL NEUROPATHY
C0041848|T047||SNOMEDCT_US|NEUROPATHY; IDIOPATHIC
C0041848|T047||SNOMEDCT_US|IDIOPATHIC NEUROPATHY
C0235024|T047|48780006|SNOMEDCT_US|NEURITIS CRANIAL|CRANIAL NEURITIS (DISORDER)
C0235024|T047|48780006|SNOMEDCT_US|CRANIAL NEURITIS|CRANIAL NEURITIS (DISORDER)
C0235024|T047|48780006|SNOMEDCT_US|CRANIAL NEURITIS |CRANIAL NEURITIS (DISORDER)
C0235024|T047|48780006|SNOMEDCT_US|CRANIAL NEURITIS, NOS|CRANIAL NEURITIS (DISORDER)
C0235880|T047|267600005|SNOMEDCT_US|MONONEURITIS OF UNSPECIFIED SITE|MONONEURITIS OF UNSPECIFIED SITE NOS (DISORDER)
C0235880|T047|267600005|SNOMEDCT_US|MONONEURITIS|MONONEURITIS OF UNSPECIFIED SITE NOS (DISORDER)
C0235880|T047|267600005|SNOMEDCT_US|MONONEURITIS |MONONEURITIS OF UNSPECIFIED SITE NOS (DISORDER)
C0235880|T047|267600005|SNOMEDCT_US|MONONEURITIDES|MONONEURITIS OF UNSPECIFIED SITE NOS (DISORDER)
C0235880|T047|267600005|SNOMEDCT_US|MONONEURITIS NOS|MONONEURITIS OF UNSPECIFIED SITE NOS (DISORDER)
C0235880|T047|267600005|SNOMEDCT_US|MONONEURITIS OF UNSPECIFIED SITE NOS |MONONEURITIS OF UNSPECIFIED SITE NOS (DISORDER)
C0235880|T047|267600005|SNOMEDCT_US|MONONEURITIS OF UNSPECIFIED SITE NOS|MONONEURITIS OF UNSPECIFIED SITE NOS (DISORDER)
C0235880|T047|267600005|SNOMEDCT_US|MONONEURITIS |MONONEURITIS OF UNSPECIFIED SITE NOS (DISORDER)
C0235880|T047|267600005|SNOMEDCT_US|MONONEURITIS, NOS|MONONEURITIS OF UNSPECIFIED SITE NOS (DISORDER)
C0270921|T047|60703000|SNOMEDCT_US|AXONAL NEUROPATHY|AXONAL NEUROPATHY (DISORDER)
C0270921|T047|60703000|SNOMEDCT_US|AXONAL NEUROPATHY |AXONAL NEUROPATHY (DISORDER)
C0270921|T047|60703000|SNOMEDCT_US|AXONAL NEUROPATHY, NOS|AXONAL NEUROPATHY (DISORDER)
C0001198|T047|66695004|SNOMEDCT_US|MERCURY POSIONING|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|FEERS DISEASE|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|SWIFTS DISEASE|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|FEERS DIS|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|SWIFTS DIS|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|PINK DIS|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|SWIFT DIS|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|FEER DIS|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|ERYTHEMA, ACRODYNIC|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|CHILDHOOD MERCURIALISM, CHRONIC|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|MERCURIALISM, CHRONIC CHILDHOOD|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|CHILDHOOD MERCURIALISMS, CHRONIC|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|CHRONIC CHILDHOOD MERCURIALISMS|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|ACRODYNIA [DISEASE/FINDING]|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|SWIFT DISEASE|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|CHRONIC CHILDHOOD MERCURIALISM|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|SWIFT'S DISEASE|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|ACRODYNIC ERYTHEMA|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|FEER'S DISEASE|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|FEER DISEASE|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|PINK DISEASE|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|SELTER'S DISEASE|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|SWIFT-FEER DISEASE|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|DISEASE PINK|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|ERYTHREDEMA POLYNEUROPATHY|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|BILDERBECK'S DISEASE|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|ACRODYNIA CAUSED BY MERCURY |ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|ACRODYNIA CAUSED BY MERCURY POISONING|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|ACRODYNIA DUE TO MERCURY |ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|ACRODYNIA DUE TO MERCURY|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|ACRODYNIA DUE TO MERCURY POISONING|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|ERYTHROEDEMA POLYNEUROPATHY|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|ACRODYNIA CAUSED BY MERCURY|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|DISEASE; PINK|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|ERYTHREDEMA; POLYNEURITIC|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|ERYTHREDEMA|ERYTHROEDEMA POLYNEUROPATHY
C0001198|T047|66695004|SNOMEDCT_US|PINK; DISEASE|ERYTHROEDEMA POLYNEUROPATHY
C0002768|T047|403605007|SNOMEDCT_US|PAIN INSENSITIVITY, CONGENITAL|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|CONGENITAL PAIN INSENSITIVITY|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|ANALGESIA CONGEN|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|PAIN INSENSITIVITY CONGEN|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|CONGEN PAIN INSENSITIVITY|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|CONGEN ANALGESIA|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|INSENSITIVITY CONGEN PAIN|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|PAIN INDIFFERENCE CONGEN|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|CONGENITAL PAIN INDIFFERENCES|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|CONGENITAL INDIFFERENCE TO PAIN|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|ANALGESIA, CONGENITAL|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|CONGENITAL ANALGESIA|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|CONGENITAL PAIN INDIFFERENCE|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|INSENSITIVITY, CONGENITAL PAIN|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|PAIN INDIFFERENCE, CONGENITAL|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|PAIN INSENSITIVITY, CONGENITAL [DISEASE/FINDING]|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|INSENSITIVITY TO PAIN, CONGENITAL|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|CHANNELOPATHY-ASSOCIATED INSENSITIVITY TO PAIN|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|CONGENITAL INSENSITIVITY TO PAIN|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|CONGENITAL INDIFFERENCE TO PAIN |CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|CONGENITAL PAIN ASYMBOLIA|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0002768|T047|403605007|SNOMEDCT_US|ASYMBOLIA|CONGENITAL INDIFFERENCE TO PAIN (FINDING)
C0027743|T047||SNOMEDCT_US|COMPRESSION SYNDROME, NERVE
C0027743|T047||SNOMEDCT_US|COMPRESSION SYNDROMES, NERVE
C0027743|T047||SNOMEDCT_US|NERVE COMPRESSION SYNDROME
C0027743|T047||SNOMEDCT_US|NERVE COMPRESSION SYNDROMES
C0027743|T047||SNOMEDCT_US|SYNDROME, NERVE COMPRESSION
C0027743|T047||SNOMEDCT_US|SYNDROMES, NERVE COMPRESSION
C0027743|T047||SNOMEDCT_US|NERVE COMPRESSION SYNDROMES [DISEASE/FINDING]
C0152025|T047|194530007|SNOMEDCT_US|POLYNEUROPATHY|[X]POLYNEUROPATHY, UNSPECIFIED (DISORDER)
C0152025|T047|194530007|SNOMEDCT_US|POLYNEUROPATHY, UNSPECIFIED|[X]POLYNEUROPATHY, UNSPECIFIED (DISORDER)
C0152025|T047|194530007|SNOMEDCT_US|POLYNEUROPATHY |[X]POLYNEUROPATHY, UNSPECIFIED (DISORDER)
C0152025|T047|194530007|SNOMEDCT_US|POLYNEUROPATHIES|[X]POLYNEUROPATHY, UNSPECIFIED (DISORDER)
C0152025|T047|194530007|SNOMEDCT_US|POLYNEUROPATHIES [DISEASE/FINDING]|[X]POLYNEUROPATHY, UNSPECIFIED (DISORDER)
C0152025|T047|194530007|SNOMEDCT_US|POLYNEUROPATHY (MULTIPLE NERVE DISORDER)|[X]POLYNEUROPATHY, UNSPECIFIED (DISORDER)
C0152025|T047|194530007|SNOMEDCT_US|POLYNEUROPATHY UNSPECIFIED|[X]POLYNEUROPATHY, UNSPECIFIED (DISORDER)
C0152025|T047|194530007|SNOMEDCT_US|POLYNEUROPATHY |[X]POLYNEUROPATHY, UNSPECIFIED (DISORDER)
C0152025|T047|194530007|SNOMEDCT_US|[X]POLYNEUROPATHY, UNSPECIFIED |[X]POLYNEUROPATHY, UNSPECIFIED (DISORDER)
C0152025|T047|194530007|SNOMEDCT_US|POLYNEUROPATHY UNSPECIFIED |[X]POLYNEUROPATHY, UNSPECIFIED (DISORDER)
C0152025|T047|194530007|SNOMEDCT_US|[X]POLYNEUROPATHY, UNSPECIFIED|[X]POLYNEUROPATHY, UNSPECIFIED (DISORDER)
C0152025|T047|194530007|SNOMEDCT_US|POLYNEUROPATHY NOS|[X]POLYNEUROPATHY, UNSPECIFIED (DISORDER)
C0152025|T047|194530007|SNOMEDCT_US|NEUROPATHY; MULTIPLE|[X]POLYNEUROPATHY, UNSPECIFIED (DISORDER)
C0152025|T047|194530007|SNOMEDCT_US|POLYNEUROPATHY, NOS|[X]POLYNEUROPATHY, UNSPECIFIED (DISORDER)
C0700594|T047|394640000|SNOMEDCT_US|RADICULOPATHY|RADICULOPATHY (DISORDER)
C0700594|T047|394640000|SNOMEDCT_US|RADICULOPATHY |RADICULOPATHY (DISORDER)
C0700594|T047|394640000|SNOMEDCT_US|RADICULOPATHIES|RADICULOPATHY (DISORDER)
C0700594|T047|394640000|SNOMEDCT_US|RADICULOPATHY, SITE UNSPECIFIED|RADICULOPATHY (DISORDER)
C0700594|T047|394640000|SNOMEDCT_US|RADICULOPATHY [DISEASE/FINDING]|RADICULOPATHY (DISORDER)
C0700594|T047|394640000|SNOMEDCT_US|RADICULAR SYNDROME|RADICULOPATHY (DISORDER)
C0700594|T047|394640000|SNOMEDCT_US|RADICULOPATHY |RADICULOPATHY (DISORDER)
C0700594|T047|394640000|SNOMEDCT_US|RADICULOPATHY NOS|RADICULOPATHY (DISORDER)
C0700594|T047|394640000|SNOMEDCT_US|SPINAL NERVE ROOT DISORDER NOS|RADICULOPATHY (DISORDER)
C0700594|T047|394640000|SNOMEDCT_US|NEUROPATHY; RADICULAR|RADICULOPATHY (DISORDER)
C0700594|T047|394640000|SNOMEDCT_US|RADICULAR; NEUROPATHIC|RADICULOPATHY (DISORDER)
C0700594|T047|394640000|SNOMEDCT_US|RADICULAR; SYNDROME|RADICULOPATHY (DISORDER)
C0700594|T047|394640000|SNOMEDCT_US|SYNDROME; RADICULAR|RADICULOPATHY (DISORDER)
C0700594|T047|394640000|SNOMEDCT_US|RADICULOPATHY, NOS|RADICULOPATHY (DISORDER)
C0206247|T047|193187004|SNOMEDCT_US|AMYLOID NEUROPATHIES|POLYNEUROPATHY IN AMYLOIDOSIS (DISORDER)
C0206247|T047|193187004|SNOMEDCT_US|AMYLOID POLYNEUROPATHY|POLYNEUROPATHY IN AMYLOIDOSIS (DISORDER)
C0206247|T047|193187004|SNOMEDCT_US|NEUROPATHY, AMYLOID|POLYNEUROPATHY IN AMYLOIDOSIS (DISORDER)
C0206247|T047|193187004|SNOMEDCT_US|POLYNEUROPATHIES, AMYLOID|POLYNEUROPATHY IN AMYLOIDOSIS (DISORDER)
C0206247|T047|193187004|SNOMEDCT_US|AMYLOID NEUROPATHY|POLYNEUROPATHY IN AMYLOIDOSIS (DISORDER)
C0206247|T047|193187004|SNOMEDCT_US|POLYNEUROPATHY, AMYLOID|POLYNEUROPATHY IN AMYLOIDOSIS (DISORDER)
C0206247|T047|193187004|SNOMEDCT_US|AMYLOID POLYNEUROPATHY |POLYNEUROPATHY IN AMYLOIDOSIS (DISORDER)
C0206247|T047|193187004|SNOMEDCT_US|AMYLOID POLYNEUROPATHIES|POLYNEUROPATHY IN AMYLOIDOSIS (DISORDER)
C0206247|T047|193187004|SNOMEDCT_US|NEUROPATHIES, AMYLOID|POLYNEUROPATHY IN AMYLOIDOSIS (DISORDER)
C0206247|T047|193187004|SNOMEDCT_US|AMYLOID NEUROPATHIES [DISEASE/FINDING]|POLYNEUROPATHY IN AMYLOIDOSIS (DISORDER)
C0206247|T047|193187004|SNOMEDCT_US|AMYLOID POLYNEUROPATHY |POLYNEUROPATHY IN AMYLOIDOSIS (DISORDER)
C0206247|T047|193187004|SNOMEDCT_US|POLYNEUROPATHY IN AMYLOIDOSIS|POLYNEUROPATHY IN AMYLOIDOSIS (DISORDER)
C0206247|T047|193187004|SNOMEDCT_US|POLYNEUROPATHY IN AMYLOIDOSIS |POLYNEUROPATHY IN AMYLOIDOSIS (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|GUILLAIN-BARRE SYNDROME|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|SYNDROME, GUILLAIN-BARRE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|GUILLAIN BARRE SYNDROME|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE IDIOPATHIC POLYNEURITIS|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|AIDP|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFLAMM POLYRADICULONEUROPATHY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|DEMYELINATING POLYRADICULONEUROPATHY ACUTE INFLAMM|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|INFLAMM POLYNEUROPATHY ACUTE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|POLYNEUROPATHY ACUTE INFLAMM|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|POLYRADICULONEUROPATHY ACUTE INFLAMM DEMYELINATING|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|INFLAMM DEMYELINATING POLYRADICULONEUROPATHY ACUTE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFLAMM POLYNEUROPATHY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|POLYRADICULONEUROPATHY ACUTE INFLAMM|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFLAMM DEMYELINATING POLYRADICULONEUROPATHY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE POSTINFECTIOUS POLYNEUROPATHY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|LANDRY'S PARALYSIS|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|POSTINFECTIOUS POLYNEURITIS|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|INFECTIOUS NEURONITIS|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFECTIOUS POLYNEURITIS |ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFECTIOUS POLYNEURITIS|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE AUTOIMMUNE NEUROPATHIES|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|AUTOIMMUNE NEUROPATHIES, ACUTE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|AUTOIMMUNE NEUROPATHY, ACUTE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|NEUROPATHIES, ACUTE AUTOIMMUNE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|NEUROPATHY, ACUTE AUTOIMMUNE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFLAMMATORY POLYNEUROPATHIES|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|INFLAMMATORY POLYNEUROPATHIES, ACUTE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|POLYNEUROPATHIES, ACUTE INFLAMMATORY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|INFLAMMATORY POLYNEUROPATHY, ACUTE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFLAMMATORY POLYRADICULONEUROPATHIES|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|INFLAMMATORY POLYRADICULONEUROPATHIES, ACUTE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|POLYRADICULONEUROPATHIES, ACUTE INFLAMMATORY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|LANDRY GUILLAIN BARRE SYNDROME|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|SYNDROME, LANDRY-GUILLAIN-BARRE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|GUILLAINE BARRE SYNDROME|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|SYNDROME, GUILLAINE-BARRE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|AC INFECT POLYNEURITIS|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE, INFLAMMATORY POLYNEUROPATHY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|POLYNEUROPATHY ACUTE, INFLAMMATORY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|INFLAMMATORY POLYNEUROPATHY ACUTES|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|INFLAMMATORY DEMYELINATING POLYRADICULONEUROPATHY, ACUTE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE AUTOIMMUNE NEUROPATHY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFLAMMATORY POLYNEUROPATHY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|DEMYELINATING POLYRADICULONEUROPATHY, ACUTE INFLAMMATORY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|POLYNEUROPATHY, ACUTE INFLAMMATORY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|POLYRADICULONEUROPATHY, ACUTE INFLAMMATORY DEMYELINATING|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|INFLAMMATORY POLYNEUROPATHY ACUTE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFLAMMATORY DEMYELINATING POLYRADICULONEUROPATHY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFLAMMATORY POLYRADICULONEUROPATHY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|POLYRADICULONEUROPATHY, ACUTE INFLAMMATORY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFLAMMATORY DEMYELINATING POLYNEUROPATHY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|INFECTIOUS POLYNEURITIS|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) |ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFECTIVE POLYNEURITIS|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INF. POLYNEURITIS|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFLAMMATORY DEMYELINATING POLYNEUROPATHY |ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFECTIVE POLYNEURITIS NOS|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFECTIVE POLYNEURITIS NOS |ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME])|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFECTIVE POLYNEURITIS |ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|POLYNEUROPATHY, INFLAMMATORY DEMYELINATING, ACUTE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFLAMMATORY DEMYELINATING POLYRADICULOPATHY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|GUILLAINE-BARRE SYNDROME|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|LANDRY-GUILLAIN-BARRE SYNDROME|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|GUILLAIN-BARRE SYNDROME, FAMILIAL|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE INFLAMMATORY NEUROPATHY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE POST-INFECTIVE RADICULONEUROPATHY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|POST-INFECTIOUS POLYNEURITIS|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|ACUTE IDIOPATHIC POLYRADICULONEURITIS|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|INFECTIOUS NEURONITIS |ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|POST-INFECTIOUS POLYNEURITIS |ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|LANDRY; PARALYSIS|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|INFECTIVE; POLYNEURITIC|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|MULTIPLE; NEURITIS, INFECTIVE, ACUTE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|NEURITIS; MULTIPLE, INFECTIVE, ACUTE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|PARALYSIS; LANDRY|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|POLYNEURITIS; ACUTE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|POLYNEURITIS; INFECTIVE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|POLYNEURITIS; POSTINFECTIVE|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|POSTINFECTIVE; POLYNEURITIC|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C3542501|T047|155082001|SNOMEDCT_US|PNS NEURONITIS|ACUTE INFECTIVE POLYNEURITIS (& [GUILLAIN-BARRE SYNDROME]) (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|ISAAC SYNDROME|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|ISAACS MERTENS SYNDROME|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|ISAACS SYNDROME|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|ISAACS-MERTENS SYNDROME|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|ISAACS SYNDROME |NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|CONTINUOUS MYOKYMIA|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|CONTINUOUS MYOKYMIAS|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|MYOKYMIAS, CONTINUOUS|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|GAMSTORP WOHLFART SYNDROME|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|ISAACS PSEUDOMYOTONIA SYNDROME|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|PSEUDOMYOTONIA|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|ISAACS SYNDROME [DISEASE/FINDING]|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|GAMSTORP-WOHLFART SYNDROME|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|ISAACS' SYNDROME|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|MYOKYMIA, CONTINUOUS|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|NEUROMYOTONIA|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|PSEUDOMYOTONIA SYNDROME OF ISAACS|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|CONTINUOUS MUSCLE ACTIVITY SYNDROME|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|SYNDROME OF CONTINUOUS MUSCLE ACTIVITY|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|QUANTAL SQUANDER|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|SYNDROMES, GAMSTORP-WOHLFART|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|SYNDROMES, ISAACS-MERTENS|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|GAMSTORP-WOHLFART SYNDROMES|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|MYOKYMIA, MYOTONIA, MUSCLE WASTING, AND HYPERHIDROSIS|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|NMAN|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|NEUROMYOTONIA AND AXONAL NEUROPATHY, AUTOSOMAL RECESSIVE|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|NEUROMYOTONIA |NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|GAMSTORP DISEASE|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|MYOKYMIA, MYOTONIA, AND MUSCLE WASTING|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|AUTOSOMAL RECESSIVE NEUROMYOTONIA WITH AXONAL NEUROPATHY|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|AUTOSOMAL RECESSIVE AXONAL NEUROPATHY WITH NEUROMYOTONIA |NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|MYOKYMIA, MYOTONIA AND MUSCLE WASTING|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|AUTOSOMAL RECESSIVE AXONAL NEUROPATHY WITH NEUROMYOTONIA|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|ISAAC'S SYNDROME|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|CONTINUOUS MUSCLE FIBER ACTIVITY|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|CONTINUOUS MUSCLE FIBRE ACTIVITY|NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|ISAACS SYNDROME |NEUROMYOTONIA (DISORDER)
C0242287|T047|305719002|SNOMEDCT_US|NEUROMYOTONIA [AMBIGUOUS]|NEUROMYOTONIA (DISORDER)
C0494491|T047|128189008|SNOMEDCT_US|MONONEUROPATHY, UNSPECIFIED|MONONEUROPATHY (DISORDER)
C0494491|T047|128189008|SNOMEDCT_US|MONONEUROPATHY|MONONEUROPATHY (DISORDER)
C0494491|T047|128189008|SNOMEDCT_US|MONONEUROPATHIES|MONONEUROPATHY (DISORDER)
C0494491|T047|128189008|SNOMEDCT_US|MONONEUROPATHIES [DISEASE/FINDING]|MONONEUROPATHY (DISORDER)
C0494491|T047|128189008|SNOMEDCT_US|MONONEUROPATHY |MONONEUROPATHY (DISORDER)
C0494491|T047|128189008|SNOMEDCT_US|MONONEUROPATHY NOS|MONONEUROPATHY (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|BRACHIAL PLEXUS NEUROPATHIES|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|BRACHIAL PLEXUS DISORDERS|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|BRACHIAL PLEXUS DIS|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|BRACHIAL PLEXUS DISEASE|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|PLEXUS DISEASE, BRACHIAL|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|PLEXUS DISEASES, BRACHIAL|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|BRACHIAL PLEXUS DISORDER|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|PLEXUS DISORDER, BRACHIAL|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|PLEXUS DISORDERS, BRACHIAL|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|BRACHIAL PLEXUS NEUROPATHY|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|NEUROPATHIES, BRACHIAL PLEXUS|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|NEUROPATHY, BRACHIAL PLEXUS|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|PLEXUS NEUROPATHIES, BRACHIAL|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|PLEXUS NEUROPATHY, BRACHIAL|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|PLEXOPATHIES, BRACHIAL|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|PLEXOPATHY, BRACHIAL|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|BRACHIAL PLEXOPATHY|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|BRACHIAL PLEXUS DISEASES|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|BRACHIAL PLEXUS NEUROPATHIES [DISEASE/FINDING]|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|BRACHIAL PLEXUS DISORDER |BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|BRACHIAL PLEXUS--DISEASES|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|BPN - BRACHIAL PLEXUS NEUROPATHY|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|BRACHIAL PLEXUS DISORDER |BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|BRACHIAL PLEXUS; NEUROPATHY|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|BRACHIAL PLEXUS; SYNDROME|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|DISEASE (OR DISORDER); PLEXUS, BRACHIAL|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|NEUROPATHY; BRACHIAL PLEXUS|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|PLEXUS BRACHIALIS; NEUROPATHIC|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|SYNDROME; BRACHIAL PLEXUS|BRACHIAL PLEXUS DISORDER (DISORDER)
C0700251|T047|3548001|SNOMEDCT_US|BRACHIAL PLEXUS NEUROPATHY, NOS|BRACHIAL PLEXUS DISORDER (DISORDER)
C0458219|T047|128200000|SNOMEDCT_US|COMPLEX REGIONAL PAIN SYNDROME NOS|COMPLEX REGIONAL PAIN SYNDROME (DISORDER)
C0458219|T047|128200000|SNOMEDCT_US|COMPLEX REGIONAL PAIN SYNDROMES|COMPLEX REGIONAL PAIN SYNDROME (DISORDER)
C0458219|T047|128200000|SNOMEDCT_US|COMPLEX REGIONAL PAIN SYNDROMES [DISEASE/FINDING]|COMPLEX REGIONAL PAIN SYNDROME (DISORDER)
C0458219|T047|128200000|SNOMEDCT_US|CRPS (COMPLEX REGIONAL PAIN SYNDROMES)|COMPLEX REGIONAL PAIN SYNDROME (DISORDER)
C0458219|T047|128200000|SNOMEDCT_US|PAIN SYNDROMES, REGIONAL COMPLEX|COMPLEX REGIONAL PAIN SYNDROME (DISORDER)
C0458219|T047|128200000|SNOMEDCT_US|CRPS|COMPLEX REGIONAL PAIN SYNDROME (DISORDER)
C0458219|T047|128200000|SNOMEDCT_US|COMPLEX REGIONAL PAIN SYNDROME|COMPLEX REGIONAL PAIN SYNDROME (DISORDER)
C0458219|T047|128200000|SNOMEDCT_US|COMPLEX REGIONAL PAIN SYNDROME (CRPS)|COMPLEX REGIONAL PAIN SYNDROME (DISORDER)
C0458219|T047|128200000|SNOMEDCT_US|COMPLEX REGIONAL PAIN SYNDROME |COMPLEX REGIONAL PAIN SYNDROME (DISORDER)
C0458219|T047|128200000|SNOMEDCT_US|COMPLEX REGIONAL PAIN SYNDROME |COMPLEX REGIONAL PAIN SYNDROME (DISORDER)
C0458219|T047|128200000|SNOMEDCT_US|COMPLEX REGIONAL PAIN SYNDROMES |COMPLEX REGIONAL PAIN SYNDROME (DISORDER)
C1363854|T047||SNOMEDCT_US|HAND ARM VIBRATION SYNDROME
C1363854|T047||SNOMEDCT_US|HAND-ARM VIBRATION SYNDROMES
C1363854|T047||SNOMEDCT_US|HAND-ARM VIBRATION SYNDROME
C1363854|T047||SNOMEDCT_US|SYNDROME, HAND-ARM VIBRATION
C1363854|T047||SNOMEDCT_US|SYNDROMES, HAND-ARM VIBRATION
C1363854|T047||SNOMEDCT_US|VIBRATION SYNDROME, HAND-ARM
C1363854|T047||SNOMEDCT_US|VIBRATION SYNDROMES, HAND-ARM
C1363854|T047||SNOMEDCT_US|HAND-ARM VIBRATION SYNDROME [DISEASE/FINDING]
C1363854|T047||SNOMEDCT_US|HAND AND ARM VIBRATION SYNDROME
C0031117|T047|42658009|SNOMEDCT_US|NERVE DISEASE, PERIPHERAL|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|NERVE DISEASES, PERIPHERAL|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NERVE DISEASE|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NERVE DISEASES|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|DISORDERS OF THE PERIPHERAL NERVOUS SYSTEM|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NERVOUS SYSTEM DISEASES|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PNS DISEASE|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NEUROPATHY|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PNS DIS|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NERVOUS SYSTEM DIS|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NERVE DIS|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PNS PERIPHERAL NERVOUS SYSTEM DIS|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NERVOUS SYSTEM DISORDER|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NEUROPATHY |DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NEUROPATHY (PHYSICAL FINDING)|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NEUROPATHIES|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|NEUROPATHY, PERIPHERAL|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|DISORDER OF PERIPHERAL NERVOUS SYSTEM NOS|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PNS DISEASES|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NERVOUS SYSTEM DISEASE|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NERVOUS SYSTEM DISEASES [DISEASE/FINDING]|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PNS (PERIPHERAL NERVOUS SYSTEM) DISEASES|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NERVOUS SYSTEM DISORDERS|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NERVE DISORDER|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PN - PERIPHERAL NEUROPATHY|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|NEUROPATHY;PERIPHERAL|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NERVE DISORDERS|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|DISORDERS OF PERIPHERAL NERVOUS SYSTEM|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|DISORDERS OF PERIPHERAL NERVOUS SYSTEM |DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NERVOUS SYSTEM DISORDERS |DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NERVOUS SYSTEM DISORDER NOS|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NERVOUS SYSTEM DISORDER NOS |DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|NERVES, PERIPHERAL--DISEASES|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|DISORDER OF PERIPHERAL NERVOUS SYSTEM|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|NEUROPATHY PERIPHERAL|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NEUROPATHY NOS|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NERVE DISORDER NOS|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM |DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NERVE DISEASE |DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|NEUROPATHY; PERIPHERAL|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL; NERVOUS SYSTEM, DISORDER|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL; NEUROPATHIC|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM, NOS|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NERVE DISORDER, NOS|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0031117|T047|42658009|SNOMEDCT_US|PERIPHERAL NEUROPATHY, NOS|DISORDER OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0852421|T047||SNOMEDCT_US|ACUTE POLYNEUROPATHY
C0852421|T047||SNOMEDCT_US|ACUTE POLYNEUROPATHIES
C0598589|T047||SNOMEDCT_US|HEREDITARY NEUROPATHY
C0598589|T047||SNOMEDCT_US|INHERITED NEUROPATHIES
C0598589|T047||SNOMEDCT_US|NEUROPATHY; HEREDITARY
C0598589|T047||SNOMEDCT_US|INHERITED NEUROPATHY
C0853004|T047||SNOMEDCT_US|PERIPHERAL NEUROPATHIES NEC
C1167650|T047||SNOMEDCT_US|POLYNEUROPATHY CHRONIC
C1167650|T047||SNOMEDCT_US|CHRONIC POLYNEUROPATHIES
C1167650|T047||SNOMEDCT_US|CHRONIC POLYNEUROPATHY
C0750944|T047|128123007|SNOMEDCT_US|PERIPHERAL AUTONOMIC NERVOUS SYSTEM DIS|DISORDER OF PERIPHERAL AUTONOMIC NERVOUS SYSTEM (DISORDER)
C0750944|T047|128123007|SNOMEDCT_US|AUTONOMIC PERIPHERAL NERVOUS SYSTEM DIS|DISORDER OF PERIPHERAL AUTONOMIC NERVOUS SYSTEM (DISORDER)
C0750944|T047|128123007|SNOMEDCT_US|AUTONOMIC PERIPHERAL NERVOUS SYSTEM DISEASES|DISORDER OF PERIPHERAL AUTONOMIC NERVOUS SYSTEM (DISORDER)
C0750944|T047|128123007|SNOMEDCT_US|DISORDER OF PERIPHERAL AUTONOMIC NERVOUS SYSTEM |DISORDER OF PERIPHERAL AUTONOMIC NERVOUS SYSTEM (DISORDER)
C0750944|T047|128123007|SNOMEDCT_US|DISORDER OF PERIPHERAL AUTONOMIC NERVOUS SYSTEM|DISORDER OF PERIPHERAL AUTONOMIC NERVOUS SYSTEM (DISORDER)
C0750944|T047|128123007|SNOMEDCT_US|DISEASE (OR DISORDER); PERIPHERAL, AUTONOMIC NERVOUS SYSTEM|DISORDER OF PERIPHERAL AUTONOMIC NERVOUS SYSTEM (DISORDER)
C0750944|T047|128123007|SNOMEDCT_US|DISORDER OF PERIPHERAL AUTONOMIC NERVOUS SYSTEM, NOS|DISORDER OF PERIPHERAL AUTONOMIC NERVOUS SYSTEM (DISORDER)
C0750944|T047|128123007|SNOMEDCT_US|PERIPHERAL AUTONOMIC NERVOUS SYSTEM DISEASES|DISORDER OF PERIPHERAL AUTONOMIC NERVOUS SYSTEM (DISORDER)
C0393912|T047|230659005|SNOMEDCT_US|AUTONOMIC DYSFUNCTION, SEGMENTAL|SEGMENTAL AUTONOMIC DYSFUNCTION (DISORDER)
C0393912|T047|230659005|SNOMEDCT_US|AUTONOMIC DYSFUNCTIONS, SEGMENTAL|SEGMENTAL AUTONOMIC DYSFUNCTION (DISORDER)
C0393912|T047|230659005|SNOMEDCT_US|SEGMENTAL AUTONOMIC DYSFUNCTIONS|SEGMENTAL AUTONOMIC DYSFUNCTION (DISORDER)
C0393912|T047|230659005|SNOMEDCT_US|SEGMENTAL AUTONOMIC DYSFUNCTION|SEGMENTAL AUTONOMIC DYSFUNCTION (DISORDER)
C0393912|T047|230659005|SNOMEDCT_US|SEGMENTAL AUTONOMIC DYSFUNCTION |SEGMENTAL AUTONOMIC DYSFUNCTION (DISORDER)
C0393918|T047|230665005|SNOMEDCT_US|DRUG-INDUCED AUTONOMIC DYSFUNCTION|DRUG-INDUCED AUTONOMIC DYSFUNCTION (DISORDER)
C0393918|T047|230665005|SNOMEDCT_US|DRUG-INDUCED AUTONOMIC DYSFUNCTION |DRUG-INDUCED AUTONOMIC DYSFUNCTION (DISORDER)
C0393920|T047|230667002|SNOMEDCT_US|CHRONIC IDIOPATHIC ANHIDROSIS|CHRONIC IDIOPATHIC ANHIDROSIS (DISORDER)
C0393920|T047|230667002|SNOMEDCT_US|CHRONIC IDIOPATHIC ANHIDROSIS |CHRONIC IDIOPATHIC ANHIDROSIS (DISORDER)
C0393921|T047|230668007|SNOMEDCT_US|IDIOPATHIC DIFFUSE HYPERHIDROSIS|IDIOPATHIC DIFFUSE HYPERHIDROSIS (DISORDER)
C0393921|T047|230668007|SNOMEDCT_US|IDIOPATHIC DIFFUSE HYPERHIDROSIS |IDIOPATHIC DIFFUSE HYPERHIDROSIS (DISORDER)
C0259749|T047|277879009|SNOMEDCT_US|AUTONOMIC NEUROPATHY|AUTONOMIC NEUROPATHY (DISORDER)
C0259749|T047|277879009|SNOMEDCT_US|AUTONOMIC NEUROPATHY NOS|AUTONOMIC NEUROPATHY (DISORDER)
C0259749|T047|277879009|SNOMEDCT_US|AUTONOMIC NEUROPATHY |AUTONOMIC NEUROPATHY (DISORDER)
C0560614|T047|282746001|SNOMEDCT_US|AUTONOMIC NERVE INJURY|AUTONOMIC NERVE INJURY (DISORDER)
C0560614|T047|282746001|SNOMEDCT_US|AUTONOMIC NERVE INJURY |AUTONOMIC NERVE INJURY (DISORDER)
C1269759|T047|371109001|SNOMEDCT_US|IMMATURE AUTONOMIC STABILITY|IMMATURE AUTONOMIC STABILITY
C1269759|T047|371109001|SNOMEDCT_US|IMMATURE AUTONOMIC SYSTEM |IMMATURE AUTONOMIC STABILITY
C1269759|T047|371109001|SNOMEDCT_US|IMMATURE AUTONOMIC SYSTEM|IMMATURE AUTONOMIC STABILITY
C0542142|T047|42998008|SNOMEDCT_US|RECURRENT LARYNGEAL NERVE PARALYSIS|VAGUS NERVE LARYNGEAL PARALYSIS (DISORDER)
C0542142|T047|42998008|SNOMEDCT_US|RECURRENT LARYNGEAL NERVE PALSY|VAGUS NERVE LARYNGEAL PARALYSIS (DISORDER)
C0542142|T047|42998008|SNOMEDCT_US|VAGUS NERVE LARYNGEAL PARALYSIS|VAGUS NERVE LARYNGEAL PARALYSIS (DISORDER)
C0542142|T047|42998008|SNOMEDCT_US|PARALYSIS RECURRENT LARYNGEAL NERVE|VAGUS NERVE LARYNGEAL PARALYSIS (DISORDER)
C0542142|T047|42998008|SNOMEDCT_US|VAGUS NERVE LARYNGEAL PARALYSIS |VAGUS NERVE LARYNGEAL PARALYSIS (DISORDER)
C0542142|T047|42998008|SNOMEDCT_US|LARYNGEAL NERVE PALSY, RECURRENT|VAGUS NERVE LARYNGEAL PARALYSIS (DISORDER)
C2317111|T047|431043000|SNOMEDCT_US|PERIPHERAL NERVE DISORDER ASSOCIATED WITH REPAIR OF HERNIA|PERIPHERAL NERVE DISORDER ASSOCIATED WITH REPAIR OF HERNIA (DISORDER)
C2317111|T047|431043000|SNOMEDCT_US|PERIPHERAL NERVE DISORDER ASSOCIATED WITH REPAIR OF HERNIA |PERIPHERAL NERVE DISORDER ASSOCIATED WITH REPAIR OF HERNIA (DISORDER)
C0393911|T047|84438001|SNOMEDCT_US|BRADBURY EGGLESTON SYNDROME|PURE AUTONOMIC FAILURE (DISORDER)
C0393911|T047|84438001|SNOMEDCT_US|SYNDROME, BRADBURY-EGGLESTON|PURE AUTONOMIC FAILURE (DISORDER)
C0393911|T047|84438001|SNOMEDCT_US|PURE AUTONOMIC FAILURE|PURE AUTONOMIC FAILURE (DISORDER)
C0393911|T047|84438001|SNOMEDCT_US|AUTONOMIC FAILURE, PURE|PURE AUTONOMIC FAILURE (DISORDER)
C0393911|T047|84438001|SNOMEDCT_US|BRADBURY-EGGLESTON SYNDROME|PURE AUTONOMIC FAILURE (DISORDER)
C0393911|T047|84438001|SNOMEDCT_US|PURE AUTONOMIC FAILURE [DISEASE/FINDING]|PURE AUTONOMIC FAILURE (DISORDER)
C0393911|T047|84438001|SNOMEDCT_US|AUTONOMIC FAILURE|PURE AUTONOMIC FAILURE (DISORDER)
C0393911|T047|84438001|SNOMEDCT_US|PURE AUTONOMIC FAILURE |PURE AUTONOMIC FAILURE (DISORDER)
C1850386|T047|128207002|SNOMEDCT_US|GIANT AXONAL NEUROPATHY 1|GIANT AXONAL NEUROPATHY (DISORDER)
C1850386|T047|128207002|SNOMEDCT_US|AXONAL NEUROPATHY, GIANT (GAN)|GIANT AXONAL NEUROPATHY (DISORDER)
C1850386|T047|128207002|SNOMEDCT_US|AXONAL NEUROPATHY, GIANT|GIANT AXONAL NEUROPATHY (DISORDER)
C1850386|T047|128207002|SNOMEDCT_US|NEUROPATHY, GIANT AXONAL (GAN)|GIANT AXONAL NEUROPATHY (DISORDER)
C1850386|T047|128207002|SNOMEDCT_US|GIANT AXONAL NEUROPATHY|GIANT AXONAL NEUROPATHY (DISORDER)
C1850386|T047|128207002|SNOMEDCT_US|GIANT AXONAL NEUROPATHY [DISEASE/FINDING]|GIANT AXONAL NEUROPATHY (DISORDER)
C1850386|T047|128207002|SNOMEDCT_US|GIANT AXONAL NEUROPATHY 1 (GAN1)|GIANT AXONAL NEUROPATHY (DISORDER)
C1850386|T047|128207002|SNOMEDCT_US|NEUROPATHY, GIANT AXONAL|GIANT AXONAL NEUROPATHY (DISORDER)
C1850386|T047|128207002|SNOMEDCT_US|GIANT AXONAL NEUROPATHY (GAN)|GIANT AXONAL NEUROPATHY (DISORDER)
C1850386|T047|128207002|SNOMEDCT_US|NEUROPATHY, GIANT AXONAL, AUTOSOMAL RECESSIVE|GIANT AXONAL NEUROPATHY (DISORDER)
C1850386|T047|128207002|SNOMEDCT_US|GIANT AXONAL NEUROPATHY 1, AUTOSOMAL RECESSIVE|GIANT AXONAL NEUROPATHY (DISORDER)
C1850386|T047|128207002|SNOMEDCT_US|GAN|GIANT AXONAL NEUROPATHY (DISORDER)
C1850386|T047|128207002|SNOMEDCT_US|GIANT AXONAL NEUROPATHY |GIANT AXONAL NEUROPATHY (DISORDER)
C1263833|T047|128193002|SNOMEDCT_US|PHRENIC NEUROPATHY|PHRENIC NERVE DISORDER (DISORDER)
C1263833|T047|128193002|SNOMEDCT_US|PHRENIC NERVE DISORDER |PHRENIC NERVE DISORDER (DISORDER)
C1263833|T047|128193002|SNOMEDCT_US|PHRENIC NERVE DISORDER|PHRENIC NERVE DISORDER (DISORDER)
C1263833|T047|128193002|SNOMEDCT_US|N.PHRENICUS; DISORDER|PHRENIC NERVE DISORDER (DISORDER)
C0338551|T047|128215004|SNOMEDCT_US|LEPROSY NEUROPATHY|LEPROSY NEUROPATHY (DISORDER)
C0338551|T047|128215004|SNOMEDCT_US|LEPROSY NEUROPATHY |LEPROSY NEUROPATHY (DISORDER)
C0542368|T047|192918007|SNOMEDCT_US|AMYLOIDOSIS WITH PERIPHERAL AUTONOMIC NEUROPATHY|AUTONOMIC NEUROPATHY DUE TO AMYLOID (DISORDER)
C0542368|T047|192918007|SNOMEDCT_US|AMYLOIDOSIS WITH PERIPHERAL AUTONOMIC NEUROPATHY |AUTONOMIC NEUROPATHY DUE TO AMYLOID (DISORDER)
C0542368|T047|192918007|SNOMEDCT_US|AUTONOMIC NEUROPATHY DUE TO AMYLOID|AUTONOMIC NEUROPATHY DUE TO AMYLOID (DISORDER)
C0542368|T047|192918007|SNOMEDCT_US|AUTONOMIC NEUROPATHY DUE TO AMYLOID |AUTONOMIC NEUROPATHY DUE TO AMYLOID (DISORDER)
C0154741|T047|155072002|SNOMEDCT_US|MONONEURITIS OF UPPER LIMB AND MONONEURITIS MULTIPLEX|MONONEURITIS OF UPPER LIMB AND MONONEURITIS MULTIPLEX (DISORDER)
C0154741|T047|155072002|SNOMEDCT_US|MONONEURITIS OF UPPER LIMB AND MONONEURITIS MULTIPLEX |MONONEURITIS OF UPPER LIMB AND MONONEURITIS MULTIPLEX (DISORDER)
C0553762|T047|193130008|SNOMEDCT_US|ANTERIOR INTEROSSEOUS NERVE SYNDROME|ANTERIOR INTEROSSEOUS NERVE LESION (DISORDER)
C0553762|T047|193130008|SNOMEDCT_US|ANTERIOR INTEROSSEOUS NERVE LESION|ANTERIOR INTEROSSEOUS NERVE LESION (DISORDER)
C0553762|T047|193130008|SNOMEDCT_US|ANTERIOR INTEROSSEOUS NERVE LESION |ANTERIOR INTEROSSEOUS NERVE LESION (DISORDER)
C0553763|T047|193139009|SNOMEDCT_US|POSTERIOR INTEROSSEOUS NERVE LESION|POSTERIOR INTEROSSEOUS NERVE LESION (DISORDER)
C0553763|T047|193139009|SNOMEDCT_US|POSTERIOR INTEROSSEOUS NERVE LESION |POSTERIOR INTEROSSEOUS NERVE LESION (DISORDER)
C0423675|T047|202796002|SNOMEDCT_US|THORACIC AND LUMBOSACRAL NEURITIS NOS |THORACIC AND LUMBOSACRAL NEURITIS (DISORDER)
C0423675|T047|202796002|SNOMEDCT_US|THORACIC AND LUMBOSACRAL NEURITIS NOS|THORACIC AND LUMBOSACRAL NEURITIS (DISORDER)
C0423675|T047|202796002|SNOMEDCT_US|THORACIC AND LUMBOSACRAL NEURITIS|THORACIC AND LUMBOSACRAL NEURITIS (DISORDER)
C0423675|T047|202796002|SNOMEDCT_US|THORACIC AND LUMBOSACRAL NEURITIS |THORACIC AND LUMBOSACRAL NEURITIS (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|INJURY TO PERIPHERAL NERVE(S) OF SHOULDER GIRDLE AND UPPER LIMB|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|INJURY TO UNSPECIFIED NERVE OF SHOULDER GIRDLE AND UPPER LIMB|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|INJURY OF NERVES AT SHOULDER AND UPPER ARM LEVEL|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|INJURY OF UNSPECIFIED NERVE AT SHOULDER AND UPPER ARM LEVEL|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|INJURY OF PERIPHERAL NERVE OF SHOULDER GIRDLE AND/OR UPPER LIMB-RETIRED|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|INJURY OF PERIPHERAL NERVE OF SHOULDER GIRDLE AND UPPER LIMB|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|INJURY OF PERIPHERAL NERVE OF SHOULDER GIRDLE AND UPPER LIMB |PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|INJURY TO UNSPECIFIED PERIPHERAL NERVE OF SHOULDER GIRDLE AND UPPER LIMB|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|INJ NERVE SHLDR/ARM NOS|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|PERIPHERAL NERVE INJURY AT SHOULDER AND UPPER ARM LEVEL |PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|PERIPHERAL NERVE INJURY AT SHOULDER AND UPPER ARM LEVEL|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|PERIPHERAL NERVE INJURY SHOULDER AND UPPER ARM LEVEL|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|SHOULDER GIRDLE PERIPHERAL NERVE INJURY|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|SHOULDER GIRDLE OR UPPER LIMB PERIPHERAL NERVE INJURY NOS|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|INJURY OF PERIPHERAL NERVE OF SHOULDER GIRDLE AND/OR UPPER LIMB |PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|INJURY OF PERIPHERAL NERVE OF SHOULDER GIRDLE AND/OR UPPER LIMB|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|ARM PERIPHERAL NERVE INJURY|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|[X]INJURY OF UNSPECIFIED NERVE AT SHOULDER AND UPPER ARM LEVEL|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM]|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|SHOULDER GIRDLE AND UPPER LIMB PERIPHERAL NERVE INJURY|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|[X]INJURY OF UNSPECIFIED NERVE AT SHOULDER AND UPPER ARM LEVEL |PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|SHOULDER GIRDLE OR UPPER LIMB PERIPHERAL NERVE INJURY NOS |PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] |PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|INJURY OF NERVES AT SHOULDER AND UPPER ARM LEVEL |PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|INJURY OF PERIPHERAL NERVE OF SHOULDER GIRDLE AND UPPER LIMB, NOS|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|INJURY TO PERIPHERAL NERVE OF SHOULDER GIRDLE AND UPPER LIMB|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0273529|T047|212252007|SNOMEDCT_US|INJURY TO PERIPHERAL NERVES OF SHOULDER GIRDLE AND UPPER LIMB|PERIPHERAL NERVE INJURY: [SHOULDER GIRDLE] &/OR [UPPER LIMB] OR [ARM] (DISORDER)
C0393802|T047|230551000|SNOMEDCT_US|HEREDITARY OR IDIOPATHIC PERIPHERAL NEUROPATHY NOS|PERIPHERAL NEUROPATHY - HEREDITARY OR IDIOPATHIC (DISORDER)
C0393802|T047|230551000|SNOMEDCT_US|PERIPHERAL NEUROPATHY - HEREDITARY OR IDIOPATHIC|PERIPHERAL NEUROPATHY - HEREDITARY OR IDIOPATHIC (DISORDER)
C0393802|T047|230551000|SNOMEDCT_US|HEREDITARY OR IDIOPATHIC PERIPHERAL NEUROPATHY NOS |PERIPHERAL NEUROPATHY - HEREDITARY OR IDIOPATHIC (DISORDER)
C0393802|T047|230551000|SNOMEDCT_US|PERIPHERAL NEUROPATHY - HEREDITARY OR IDIOPATHIC |PERIPHERAL NEUROPATHY - HEREDITARY OR IDIOPATHIC (DISORDER)
C2239188|T047|230570005|SNOMEDCT_US|BURNING, FEET SYNDROME|BURNING FEET SYNDROME (DISORDER)
C2239188|T047|230570005|SNOMEDCT_US|BURNING FEET SYNDROME|BURNING FEET SYNDROME (DISORDER)
C2239188|T047|230570005|SNOMEDCT_US|BURNING FEET SYNDROME |BURNING FEET SYNDROME (DISORDER)
C2239188|T047|230570005|SNOMEDCT_US|STRACHAN'S SYNDROME|BURNING FEET SYNDROME (DISORDER)
C2239188|T047|230570005|SNOMEDCT_US|BURNING FEET; SYNDROME|BURNING FEET SYNDROME (DISORDER)
C2239188|T047|230570005|SNOMEDCT_US|BURNING; FEET SYNDROME|BURNING FEET SYNDROME (DISORDER)
C2239188|T047|230570005|SNOMEDCT_US|FOOT; BURNING |BURNING FEET SYNDROME (DISORDER)
C2239188|T047|230570005|SNOMEDCT_US|FOOT; SYNDROME, BURNING|BURNING FEET SYNDROME (DISORDER)
C2239188|T047|230570005|SNOMEDCT_US|SYNDROME; BURNING FEET|BURNING FEET SYNDROME (DISORDER)
C0338553|T047|230597003|SNOMEDCT_US|INTERCOSTAL POST-HERPETIC NEURALGIA|INTERCOSTAL POST-HERPETIC NEURALGIA (DISORDER)
C0338553|T047|230597003|SNOMEDCT_US|INTERCOSTAL POST-HERPETIC NEURALGIA |INTERCOSTAL POST-HERPETIC NEURALGIA (DISORDER)
C0472363|T047|230606008|SNOMEDCT_US|ISCHAEMIC NEUROPATHY DUE TO ARTERIAL STEAL|ISCHEMIC NEUROPATHY DUE TO ARTERIAL STEAL (DISORDER)
C0472363|T047|230606008|SNOMEDCT_US|ISCHEMIC NEUROPATHY DUE TO ARTERIAL STEAL|ISCHEMIC NEUROPATHY DUE TO ARTERIAL STEAL (DISORDER)
C0472363|T047|230606008|SNOMEDCT_US|ISCHEMIC NEUROPATHY DUE TO ARTERIAL STEAL |ISCHEMIC NEUROPATHY DUE TO ARTERIAL STEAL (DISORDER)
C0553760|T047|230617009|SNOMEDCT_US|LUMBOSACRAL PLEXUS NEUROPATHY|LUMBOSACRAL PLEXUS NEUROPATHY (DISORDER)
C0553760|T047|230617009|SNOMEDCT_US|LUMBOSACRAL PLEXUS NEUROPATHY |LUMBOSACRAL PLEXUS NEUROPATHY (DISORDER)
C0393880|T047|230627003|SNOMEDCT_US|PERIPHERAL NERVE COMPRESSION ARM|COMPRESSION NEUROPATHY OF UPPER LIMB (DISORDER)
C0393880|T047|230627003|SNOMEDCT_US|COMPRESSION NEUROPATHY OF UPPER LIMB|COMPRESSION NEUROPATHY OF UPPER LIMB (DISORDER)
C0393880|T047|230627003|SNOMEDCT_US|COMPRESSION NEUROPATHY OF UPPER LIMB |COMPRESSION NEUROPATHY OF UPPER LIMB (DISORDER)
C0393896|T047|230645003|SNOMEDCT_US|COMPRESSION NEUROPATHY OF TRUNK|COMPRESSION NEUROPATHY OF TRUNK (DISORDER)
C0393896|T047|230645003|SNOMEDCT_US|COMPRESSION NEUROPATHY OF TRUNK |COMPRESSION NEUROPATHY OF TRUNK (DISORDER)
C0393897|T047|230646002|SNOMEDCT_US|INTERCOSTAL NEUROPATHY|INTERCOSTAL NEUROPATHY (DISORDER)
C0393897|T047|230646002|SNOMEDCT_US|INTERCOSTAL NEUROPATHY |INTERCOSTAL NEUROPATHY (DISORDER)
C0393897|T047|230646002|SNOMEDCT_US|INTERCOSTAL NEUROPATHY |INTERCOSTAL NEUROPATHY (DISORDER)
C0393897|T047|230646002|SNOMEDCT_US|DISEASE (OR DISORDER); INTERCOSTAL NERVE|INTERCOSTAL NEUROPATHY (DISORDER)
C0393919|T047|230666006|SNOMEDCT_US|PARANEOPL AUTONOMIC DYSFUNCTION|PARANEOPLASTIC AUTONOMIC DYSFUNCTION (DISORDER)
C0393919|T047|230666006|SNOMEDCT_US|AUTONOMIC DYSFUNCTION PARANEOPL|PARANEOPLASTIC AUTONOMIC DYSFUNCTION (DISORDER)
C0393919|T047|230666006|SNOMEDCT_US|AUTONOMIC DYSFUNCTIONS, PARANEOPLASTIC|PARANEOPLASTIC AUTONOMIC DYSFUNCTION (DISORDER)
C0393919|T047|230666006|SNOMEDCT_US|PARANEOPLASTIC AUTONOMIC DYSFUNCTIONS|PARANEOPLASTIC AUTONOMIC DYSFUNCTION (DISORDER)
C0393919|T047|230666006|SNOMEDCT_US|AUTONOMIC DYSFUNCTION, PARANEOPLASTIC|PARANEOPLASTIC AUTONOMIC DYSFUNCTION (DISORDER)
C0393919|T047|230666006|SNOMEDCT_US|PARANEOPLASTIC AUTONOMIC DYSFUNCTION|PARANEOPLASTIC AUTONOMIC DYSFUNCTION (DISORDER)
C0393919|T047|230666006|SNOMEDCT_US|PARANEOPLASTIC AUTONOMIC DYSFUNCTION |PARANEOPLASTIC AUTONOMIC DYSFUNCTION (DISORDER)
C0270922|T047|23414001|SNOMEDCT_US|DEMYELINATING PERIPHERAL NEUROPATHY|PERIPHERAL DEMYELINATING NEUROPATHY (DISORDER)
C0270922|T047|23414001|SNOMEDCT_US|DEMYELINATING NEUROPATHY|PERIPHERAL DEMYELINATING NEUROPATHY (DISORDER)
C0270922|T047|23414001|SNOMEDCT_US|PERIPHERAL DEMYELINATING NEUROPATHY|PERIPHERAL DEMYELINATING NEUROPATHY (DISORDER)
C0270922|T047|23414001|SNOMEDCT_US|DEMYELINATING POLYNEUROPATHY|PERIPHERAL DEMYELINATING NEUROPATHY (DISORDER)
C0270922|T047|23414001|SNOMEDCT_US|DEMYELINATING POLYNEUROPATHY NOS|PERIPHERAL DEMYELINATING NEUROPATHY (DISORDER)
C0270922|T047|23414001|SNOMEDCT_US|PERIPHERAL DEMYELINATING NEUROPATHY |PERIPHERAL DEMYELINATING NEUROPATHY (DISORDER)
C0270922|T047|23414001|SNOMEDCT_US|DEMYELINATING NEUROPATHY, NOS|PERIPHERAL DEMYELINATING NEUROPATHY (DISORDER)
C0270922|T047|23414001|SNOMEDCT_US|DEMYELINATING POLYNEUROPATHY, NOS|PERIPHERAL DEMYELINATING NEUROPATHY (DISORDER)
C0266517|T047|23880008|SNOMEDCT_US|CONGENITAL PERIPHERAL NERVE DISORDERS|CONGENITAL ANOMALY OF PERIPHERAL NERVE (DISORDER)
C0266517|T047|23880008|SNOMEDCT_US|CONGENITAL ANOMALY OF PERIPHERAL NERVE |CONGENITAL ANOMALY OF PERIPHERAL NERVE (DISORDER)
C0266517|T047|23880008|SNOMEDCT_US|CONGENITAL ANOMALY OF PERIPHERAL NERVE|CONGENITAL ANOMALY OF PERIPHERAL NERVE (DISORDER)
C0266517|T047|23880008|SNOMEDCT_US|CONGENITAL ANOMALY OF NERVE, NOS|CONGENITAL ANOMALY OF PERIPHERAL NERVE (DISORDER)
C0413275|T047|241996007|SNOMEDCT_US|PERIPHERAL NERVE DECOMPRESSION INJURY|PERIPHERAL NERVE DECOMPRESSION INJURY (DISORDER)
C0413275|T047|241996007|SNOMEDCT_US|PERIPHERAL NERVE DECOMPRESSION INJURY |PERIPHERAL NERVE DECOMPRESSION INJURY (DISORDER)
C0423709|T047|247387008|SNOMEDCT_US|CRURALGIA|CRURALGIA (DISORDER)
C0423709|T047|247387008|SNOMEDCT_US|CRURALGIA |CRURALGIA (DISORDER)
C0344306|T047|247389006|SNOMEDCT_US|INTERCOSTAL NEURALGIA|INTERCOSTAL NEURALGIA (DISORDER)
C0344306|T047|247389006|SNOMEDCT_US|INTERCOSTAL NEURALGIA |INTERCOSTAL NEURALGIA (DISORDER)
C0394021|T047|271971004|SNOMEDCT_US|DISORDER OF PERIPHERAL NERVE GRAFT|DISORDER OF PERIPHERAL NERVE GRAFT (DISORDER)
C0394021|T047|271971004|SNOMEDCT_US|DISORDER OF PERIPHERAL NERVE GRAFT |DISORDER OF PERIPHERAL NERVE GRAFT (DISORDER)
C0565585|T047|288234009|SNOMEDCT_US|NEURALGIA/NEURITIS - SHOULDER |NEURALGIA/NEURITIS - SHOULDER (DISORDER)
C0565585|T047|288234009|SNOMEDCT_US|NEURALGIA/NEURITIS - SHOULDER|NEURALGIA/NEURITIS - SHOULDER (DISORDER)
C0565586|T047|288235005|SNOMEDCT_US|NEURALGIA/NEURITIS - UPPER ARM |NEURALGIA/NEURITIS - UPPER ARM (DISORDER)
C0565586|T047|288235005|SNOMEDCT_US|NEURALGIA/NEURITIS - UPPER ARM|NEURALGIA/NEURITIS - UPPER ARM (DISORDER)
C0565590|T047|288239004|SNOMEDCT_US|NEURALGIA/NEURITIS - LOWER LEG|NEURALGIA/NEURITIS - LOWER LEG (DISORDER)
C0565590|T047|288239004|SNOMEDCT_US|NEURALGIA/NEURITIS - LOWER LEG |NEURALGIA/NEURITIS - LOWER LEG (DISORDER)
C0565591|T047|288240002|SNOMEDCT_US|NEURALGIA/NEURITIS -ANKLE/FOOT|NEURALGIA/NEURITIS - ANKLE/FOOT (DISORDER)
C0565591|T047|288240002|SNOMEDCT_US|NEURALGIA/NEURITIS - ANKLE/FOOT|NEURALGIA/NEURITIS - ANKLE/FOOT (DISORDER)
C0565591|T047|288240002|SNOMEDCT_US|NEURALGIA/NEURITIS - ANKLE/FOOT |NEURALGIA/NEURITIS - ANKLE/FOOT (DISORDER)
C0574717|T047|297945000|SNOMEDCT_US|UPPER LIMB NERVE LESION|UPPER LIMB NERVE LESION (DISORDER)
C0574717|T047|297945000|SNOMEDCT_US|UPPER LIMB NERVE LESION |UPPER LIMB NERVE LESION (DISORDER)
C0574718|T047|297946004|SNOMEDCT_US|LOWER LIMB NERVE LESION|LOWER LIMB NERVE LESION (DISORDER)
C0574718|T047|297946004|SNOMEDCT_US|LOWER LIMB NERVE LESION |LOWER LIMB NERVE LESION (DISORDER)
C0574920|T047|298137008|SNOMEDCT_US|THORACOABDOMINAL NEUROPATHY|THORACOABDOMINAL NEUROPATHY (DISORDER)
C0574920|T047|298137008|SNOMEDCT_US|THORACOABDOMINAL NEUROPATHY |THORACOABDOMINAL NEUROPATHY (DISORDER)
C0153097|T047|31524007|SNOMEDCT_US|POLYNEUROPATHY DUE TO MUMPS|MUMPS POLYNEUROPATHY (DISORDER)
C0153097|T047|31524007|SNOMEDCT_US|POLYNEUROPATHY DUE TO MUMPS |MUMPS POLYNEUROPATHY (DISORDER)
C0153097|T047|31524007|SNOMEDCT_US|POLYNEUROPATHY MUMPS|MUMPS POLYNEUROPATHY (DISORDER)
C0153097|T047|31524007|SNOMEDCT_US|MUMPS POLYNEUROPATHY|MUMPS POLYNEUROPATHY (DISORDER)
C0153097|T047|31524007|SNOMEDCT_US|POLYNEUROPATHY IN MUMPS |MUMPS POLYNEUROPATHY (DISORDER)
C0153097|T047|31524007|SNOMEDCT_US|POLYNEUROPATHY IN MUMPS|MUMPS POLYNEUROPATHY (DISORDER)
C0153097|T047|31524007|SNOMEDCT_US|MUMPS POLYNEUROPATHY |MUMPS POLYNEUROPATHY (DISORDER)
C0271686|T047|50620007|SNOMEDCT_US|DIABETIC AUTONOMIC NEUROPATHY|DIABETIC AUTONOMIC NEUROPATHY (DISORDER)
C0271686|T047|50620007|SNOMEDCT_US|DIABETES MELLITUS WITH AUTONOMIC NEUROPATHY |DIABETIC AUTONOMIC NEUROPATHY (DISORDER)
C0271686|T047|50620007|SNOMEDCT_US|DIABETES MELLITUS WITH AUTONOMIC NEUROPATHY|DIABETIC AUTONOMIC NEUROPATHY (DISORDER)
C0271686|T047|50620007|SNOMEDCT_US|AUTONOMIC NEUROPATHIES, DIABETIC|DIABETIC AUTONOMIC NEUROPATHY (DISORDER)
C0271686|T047|50620007|SNOMEDCT_US|AUTONOMIC NEUROPATHY, DIABETIC|DIABETIC AUTONOMIC NEUROPATHY (DISORDER)
C0271686|T047|50620007|SNOMEDCT_US|DIABETIC AUTONOMIC NEUROPATHIES|DIABETIC AUTONOMIC NEUROPATHY (DISORDER)
C0271686|T047|50620007|SNOMEDCT_US|NEUROPATHIES, DIABETIC AUTONOMIC|DIABETIC AUTONOMIC NEUROPATHY (DISORDER)
C0271686|T047|50620007|SNOMEDCT_US|NEUROPATHY, DIABETIC AUTONOMIC|DIABETIC AUTONOMIC NEUROPATHY (DISORDER)
C0271686|T047|50620007|SNOMEDCT_US|AUTONOMIC NEUROPATHY DUE TO DIABETES|DIABETIC AUTONOMIC NEUROPATHY (DISORDER)
C0271686|T047|50620007|SNOMEDCT_US|DIABETIC AUTONOMIC NEUROPATHY |DIABETIC AUTONOMIC NEUROPATHY (DISORDER)
C0037887|T047|61830005|SNOMEDCT_US|SPHENOPALATINE NEURALGIA|SPHENOPALATINE NEURALGIA (DISORDER)
C0037887|T047|61830005|SNOMEDCT_US|NEURALGIA, SPHENOPALATINE|SPHENOPALATINE NEURALGIA (DISORDER)
C0037887|T047|61830005|SNOMEDCT_US|NEURALGIAS, SPHENOPALATINE|SPHENOPALATINE NEURALGIA (DISORDER)
C0037887|T047|61830005|SNOMEDCT_US|SPHENOPALATINE NEURALGIAS|SPHENOPALATINE NEURALGIA (DISORDER)
C0037887|T047|61830005|SNOMEDCT_US|SLUDER'S NEURALGIA|SPHENOPALATINE NEURALGIA (DISORDER)
C0037887|T047|61830005|SNOMEDCT_US|SPHENOPALATINE GANGLION NEURALGIA|SPHENOPALATINE NEURALGIA (DISORDER)
C0037887|T047|61830005|SNOMEDCT_US|SLUDER'S SYNDROME|SPHENOPALATINE NEURALGIA (DISORDER)
C0037887|T047|61830005|SNOMEDCT_US|SPHENOPALATINE NEURALGIA |SPHENOPALATINE NEURALGIA (DISORDER)
C0037887|T047|61830005|SNOMEDCT_US|NEURALGIA; SPHENOPALATINE|SPHENOPALATINE NEURALGIA (DISORDER)
C0037887|T047|61830005|SNOMEDCT_US|SPHENOPALATINE; NEURALGIA|SPHENOPALATINE NEURALGIA (DISORDER)
C1527351|T047|72274001|SNOMEDCT_US|NERVE ROOT DIS|NERVE ROOT DISORDER (DISORDER)
C1527351|T047|72274001|SNOMEDCT_US|NERVE ROOT DISORDERS|NERVE ROOT DISORDER (DISORDER)
C1527351|T047|72274001|SNOMEDCT_US|NERVE ROOT DISORDER|NERVE ROOT DISORDER (DISORDER)
C1527351|T047|72274001|SNOMEDCT_US|NERVE ROOT DISORDER |NERVE ROOT DISORDER (DISORDER)
C1527351|T047|72274001|SNOMEDCT_US|NERVE ROOT DISORDER, NOS|NERVE ROOT DISORDER (DISORDER)
C0262593|T047|73590005|SNOMEDCT_US|PERIPHERAL NERVE INJURY|PERIPHERAL NERVE INJURY (DISORDER)
C0262593|T047|73590005|SNOMEDCT_US|INJURY OF PERIPHERAL NERVE |PERIPHERAL NERVE INJURY (DISORDER)
C0262593|T047|73590005|SNOMEDCT_US|INJURY OF PERIPHERAL NERVE|PERIPHERAL NERVE INJURY (DISORDER)
C0262593|T047|73590005|SNOMEDCT_US|INJURY;NERVE;PERIPHERAL|PERIPHERAL NERVE INJURY (DISORDER)
C0262593|T047|73590005|SNOMEDCT_US|NERVE INJURIES, PERIPHERAL|PERIPHERAL NERVE INJURY (DISORDER)
C0262593|T047|73590005|SNOMEDCT_US|NERVE INJURY, PERIPHERAL|PERIPHERAL NERVE INJURY (DISORDER)
C0262593|T047|73590005|SNOMEDCT_US|INJURY, PERIPHERAL NERVE|PERIPHERAL NERVE INJURY (DISORDER)
C0262593|T047|73590005|SNOMEDCT_US|INJURIES, PERIPHERAL NERVE|PERIPHERAL NERVE INJURY (DISORDER)
C0262593|T047|73590005|SNOMEDCT_US|PERIPHERAL NERVE INJURIES|PERIPHERAL NERVE INJURY (DISORDER)
C0262593|T047|73590005|SNOMEDCT_US|PERIPHERAL NERVE INJURIES [DISEASE/FINDING]|PERIPHERAL NERVE INJURY (DISORDER)
C0262593|T047|73590005|SNOMEDCT_US|PERIPHERAL NERVE INJURY NOS|PERIPHERAL NERVE INJURY (DISORDER)
C0262593|T047|73590005|SNOMEDCT_US|PERIPHERAL NERVE INJURY NOS |PERIPHERAL NERVE INJURY (DISORDER)
C0262593|T047|73590005|SNOMEDCT_US|PERIPHERAL NERVE INJURY |PERIPHERAL NERVE INJURY (DISORDER)
C0262593|T047|73590005|SNOMEDCT_US|PNI - PERIPHERAL NERVE INJURY|PERIPHERAL NERVE INJURY (DISORDER)
C0262593|T047|73590005|SNOMEDCT_US|INJURY; NERVE, PERIPHERAL|PERIPHERAL NERVE INJURY (DISORDER)
C0262593|T047|73590005|SNOMEDCT_US|NERVE; INJURY, PERIPHERAL|PERIPHERAL NERVE INJURY (DISORDER)
C0262593|T047|73590005|SNOMEDCT_US|PERIPHERAL NERVE INJURY, NOS|PERIPHERAL NERVE INJURY (DISORDER)
C0338536|T047|95669001|SNOMEDCT_US|NEURALGIA SUPERIOR LARYNGEAL|SUPERIOR LARYNGEAL NEURALGIA (DISORDER)
C0338536|T047|95669001|SNOMEDCT_US|SUPERIOR LARYNGEAL NEURALGIA |SUPERIOR LARYNGEAL NEURALGIA (DISORDER)
C0338536|T047|95669001|SNOMEDCT_US|SUPERIOR LARYNGEAL NEURALGIA|SUPERIOR LARYNGEAL NEURALGIA (DISORDER)
C0338536|T047|95669001|SNOMEDCT_US|SUPERIOR LARYNGEAL NEURALGIA |SUPERIOR LARYNGEAL NEURALGIA (DISORDER)
C0270910|T047|22722001|SNOMEDCT_US|IDIOPATHIC PERIPHERAL NEUROPATHY|IDIOPATHIC PERIPHERAL NEUROPATHY (DISORDER)
C0270910|T047|22722001|SNOMEDCT_US|IDIOPATHIC PERIPHERAL NEUROPATHY |IDIOPATHIC PERIPHERAL NEUROPATHY (DISORDER)
C0270910|T047|22722001|SNOMEDCT_US|IDIOPATHIC PERIPHERAL NEUROPATHY |IDIOPATHIC PERIPHERAL NEUROPATHY (DISORDER)
C0270910|T047|22722001|SNOMEDCT_US|NEUROPATHY; PERIPHERAL, IDIOPATHIC|IDIOPATHIC PERIPHERAL NEUROPATHY (DISORDER)
C0270910|T047|22722001|SNOMEDCT_US|IDIOPATHIC PERIPHERAL NEUROPATHY, NOS|IDIOPATHIC PERIPHERAL NEUROPATHY (DISORDER)
C0795950|T047|702439002|SNOMEDCT_US|AGENESIS OF THE CORPUS CALLOSUM WITH PERIPHERAL NEUROPATHY|AGENESIS OF CORPUS CALLOSUM WITH PERIPHERAL NEUROPATHY
C0795950|T047|702439002|SNOMEDCT_US|CORPUS CALLOSUM AGENESIS NEURONOPATHY|AGENESIS OF CORPUS CALLOSUM WITH PERIPHERAL NEUROPATHY
C0795950|T047|702439002|SNOMEDCT_US|ANDERMANN SYNDROME|AGENESIS OF CORPUS CALLOSUM WITH PERIPHERAL NEUROPATHY
C0795950|T047|702439002|SNOMEDCT_US|CHARLEVOIX DISEASE|AGENESIS OF CORPUS CALLOSUM WITH PERIPHERAL NEUROPATHY
C0795950|T047|702439002|SNOMEDCT_US|POLYNEUROPATHY, SENSORIMOTOR, WITH OR WITHOUT AGENESIS OF THE CORPUS CALLOSUM|AGENESIS OF CORPUS CALLOSUM WITH PERIPHERAL NEUROPATHY
C0795950|T047|702439002|SNOMEDCT_US|CORPUS CALLOSUM, AGENESIS OF, WITH NEURONOPATHY|AGENESIS OF CORPUS CALLOSUM WITH PERIPHERAL NEUROPATHY
C0795950|T047|702439002|SNOMEDCT_US|AGENESIS OF CORPUS CALLOSUM WITH PERIPHERAL NEUROPATHY|AGENESIS OF CORPUS CALLOSUM WITH PERIPHERAL NEUROPATHY
C0795950|T047|702439002|SNOMEDCT_US|AGENESIS OF CORPUS CALLOSUM WITH POLYNEUROPATHY|AGENESIS OF CORPUS CALLOSUM WITH PERIPHERAL NEUROPATHY
C0795950|T047|702439002|SNOMEDCT_US|AGENESIS OF CORPUS CALLOSUM WITH NEURONOPATHY|AGENESIS OF CORPUS CALLOSUM WITH PERIPHERAL NEUROPATHY
C0795950|T047|702439002|SNOMEDCT_US|HEREDITARY MOTOR AND SENSORY NEUROPATHY WITH AGENESIS OF THE CORPUS CALLOSUM|AGENESIS OF CORPUS CALLOSUM WITH PERIPHERAL NEUROPATHY
C0795950|T047|702439002|SNOMEDCT_US|AGENESIS OF CORPUS CALLOSUM WITH PERIPHERAL NEUROPATHY |AGENESIS OF CORPUS CALLOSUM WITH PERIPHERAL NEUROPATHY
C0796123|T047||SNOMEDCT_US|CATARACT-ATAXIA-DEAFNESS-RETARDATION SYNDROME
C0796123|T047||SNOMEDCT_US|CATARACT ATAXIA DEAFNESS
C0796123|T047||SNOMEDCT_US|BEGEER SYNDROME
C0796123|T047||SNOMEDCT_US|CATARACT ATAXIA DEAFNESS SYNDROME
C0796123|T047||SNOMEDCT_US|POLYNEUROPATHY, CATARACT, DEAFNESS SYNDROME
C0796123|T047||SNOMEDCT_US|POLYNEUROPATHY-CATARACT-DEAFNESS SYNDROME
C1850406|T047||SNOMEDCT_US|NAVAJO NEUROHEPATOPATHY
C1850406|T047||SNOMEDCT_US|NAVAJO NEUROPATHY
C1850406|T047||SNOMEDCT_US|MITOCHONDRIAL DNA DEPLETION SYNDROME 6 (HEPATOCEREBRAL TYPE)
C1850406|T047||SNOMEDCT_US|MTDPS6
C1850406|T047||SNOMEDCT_US|MPV17-ASSOCIATED HEPATOCEREBRAL MDS
C1850406|T047||SNOMEDCT_US|MPV17-RELATED HEPATOCEREBRAL MITOCHONDRIAL DNA DEPLETION SYNDROME
C1850406|T047||SNOMEDCT_US|MITOCHONDRIAL DNA DEPLETION SYNDROME 6
C2932678|T047||SNOMEDCT_US|INHERITED PERIPHERAL NEUROPATHY
C0006091|T047|193109004|SNOMEDCT_US|BRACHIAL PLEXUS LESIONS|BRACHIAL PLEXUS LESIONS NOS (DISORDER)
C0006091|T047|193109004|SNOMEDCT_US|LESION;BRACHIAL PLEXUS|BRACHIAL PLEXUS LESIONS NOS (DISORDER)
C0006091|T047|193109004|SNOMEDCT_US|BRACHIAL PLEXUS LESIONS NOS|BRACHIAL PLEXUS LESIONS NOS (DISORDER)
C0006091|T047|193109004|SNOMEDCT_US|BRACHIAL PLEXUS LESIONS NOS |BRACHIAL PLEXUS LESIONS NOS (DISORDER)
C0006091|T047|193109004|SNOMEDCT_US|BRACHIAL PLEXUS LESION|BRACHIAL PLEXUS LESIONS NOS (DISORDER)
C0006091|T047|193109004|SNOMEDCT_US|BRACHIAL PLEXUS; LESION|BRACHIAL PLEXUS LESIONS NOS (DISORDER)
C0006091|T047|193109004|SNOMEDCT_US|LESION; BRACHIAL PLEXUS|BRACHIAL PLEXUS LESIONS NOS (DISORDER)
C0006091|T047|193109004|SNOMEDCT_US|PLEXUS BRACHIALIS; LESION|BRACHIAL PLEXUS LESIONS NOS (DISORDER)
C0006091|T047|193109004|SNOMEDCT_US|BRACHIAL PLEXUS LESION, NOS|BRACHIAL PLEXUS LESIONS NOS (DISORDER)
C0006091|T047|193109004|SNOMEDCT_US|LESION OF BRACHIAL PLEXUS|BRACHIAL PLEXUS LESIONS NOS (DISORDER)
C2959948|T047|446494003|SNOMEDCT_US|EPENDYMAL CYST OF SPINAL NERVE |EPENDYMAL CYST OF SPINAL NERVE (DISORDER)
C2959948|T047|446494003|SNOMEDCT_US|EPENDYMAL CYST OF SPINAL NERVE|EPENDYMAL CYST OF SPINAL NERVE (DISORDER)
C0271676|T047|78409004|SNOMEDCT_US|ABDOMINAL POLYRADICULOPATHIES|ABDOMINAL POLYRADICULOPATHY (DISORDER)
C0271676|T047|78409004|SNOMEDCT_US|ABDOMINAL POLYRADICULOPATHY|ABDOMINAL POLYRADICULOPATHY (DISORDER)
C0271676|T047|78409004|SNOMEDCT_US|POLYRADICULOPATHIES, ABDOMINAL|ABDOMINAL POLYRADICULOPATHY (DISORDER)
C0271676|T047|78409004|SNOMEDCT_US|ABDOMINAL POLYRADICULOPATHY |ABDOMINAL POLYRADICULOPATHY (DISORDER)
C0271676|T047|78409004|SNOMEDCT_US|POLYRADICULOPATHY, ABDOMINAL|ABDOMINAL POLYRADICULOPATHY (DISORDER)
C2119284|T047||SNOMEDCT_US|UNCONTROLLED TYPE I DIABETES MELLITUS WITH PERIPHERAL NEUROPATHY 
C2119284|T047||SNOMEDCT_US|TYPE 1 DIABETIC PERIPHERAL NEUROPATHY, UNCONTROLLED
C2119284|T047||SNOMEDCT_US|UNCONTROLLED TYPE 1 DIABETES MELLITUS WITH PERIPHERAL NEUROPATHY 
C2119284|T047||SNOMEDCT_US|UNCONTROLLED TYPE 1 DIABETES MELLITUS WITH PERIPHERAL NEUROPATHY
C1827029|T047|423023005|SNOMEDCT_US|ENTRAPMENT NEUROPATHY OF UPPER LIMB |ENTRAPMENT NEUROPATHY OF UPPER LIMB (DISORDER)
C1827029|T047|423023005|SNOMEDCT_US|ENTRAPMENT NEUROPATHY OF UPPER LIMB|ENTRAPMENT NEUROPATHY OF UPPER LIMB (DISORDER)
C0154758|T047|267601009|SNOMEDCT_US|INFLAMMATORY AND TOXIC NEUROPATHY|INFLAMMATORY AND TOXIC NEUROPATHY (DISORDER)
C0154758|T047|267601009|SNOMEDCT_US|UNSPECIFIED INFLAMMATORY AND TOXIC NEUROPATHIES|INFLAMMATORY AND TOXIC NEUROPATHY (DISORDER)
C0154758|T047|267601009|SNOMEDCT_US|INFLAM/TOX NEUROPTHY NOS|INFLAMMATORY AND TOXIC NEUROPATHY (DISORDER)
C0154758|T047|267601009|SNOMEDCT_US|UNSPECIFIED INFLAMMATORY AND TOXIC NEUROPATHY|INFLAMMATORY AND TOXIC NEUROPATHY (DISORDER)
C0154758|T047|267601009|SNOMEDCT_US|INFLAMMATORY &/OR TOXIC NEUROPATHY |INFLAMMATORY AND TOXIC NEUROPATHY (DISORDER)
C0154758|T047|267601009|SNOMEDCT_US|TOXIC OR INFLAMMATORY NEUROPATHY NOS|INFLAMMATORY AND TOXIC NEUROPATHY (DISORDER)
C0154758|T047|267601009|SNOMEDCT_US|TOXIC OR INFLAMMATORY NEUROPATHY NOS |INFLAMMATORY AND TOXIC NEUROPATHY (DISORDER)
C0154758|T047|267601009|SNOMEDCT_US|INFLAMMATORY &/OR TOXIC NEUROPATHY|INFLAMMATORY AND TOXIC NEUROPATHY (DISORDER)
C0154758|T047|267601009|SNOMEDCT_US|INFLAMMATORY AND TOXIC NEUROPATHY |INFLAMMATORY AND TOXIC NEUROPATHY (DISORDER)
C0270109|T047|28778005|SNOMEDCT_US|PHRENIC NERVE PARALYSIS DUE TO BIRTH INJURY|PHRENIC NERVE PARALYSIS AS BIRTH TRAUMA (DISORDER)
C0270109|T047|28778005|SNOMEDCT_US|PHRENIC NERVE PARALYSIS AS BIRTH TRAUMA|PHRENIC NERVE PARALYSIS AS BIRTH TRAUMA (DISORDER)
C0270109|T047|28778005|SNOMEDCT_US|PHRENIC NERVE PARALYSIS AS BIRTH TRAUMA |PHRENIC NERVE PARALYSIS AS BIRTH TRAUMA (DISORDER)
C0270109|T047|28778005|SNOMEDCT_US|PHRENIC NERVE PARALYSIS DUE TO BIRTH TRAUMA|PHRENIC NERVE PARALYSIS AS BIRTH TRAUMA (DISORDER)
C0393852|T047|230595006|SNOMEDCT_US|NEUROPATHY DUE TO INFECTION|NEUROPATHY DUE TO INFECTION (DISORDER)
C0393852|T047|230595006|SNOMEDCT_US|NEUROPATHY DUE TO INFECTION |NEUROPATHY DUE TO INFECTION (DISORDER)
C0273522|T047|212191006|SNOMEDCT_US|CAUDA EQUINA INJURY WITHOUT BONY INJURY |CAUDA EQUINA INJURY WITHOUT BONY INJURY (DISORDER)
C0273522|T047|212191006|SNOMEDCT_US|CAUDA EQUINA INJURY WITHOUT BONY INJURY|CAUDA EQUINA INJURY WITHOUT BONY INJURY (DISORDER)
C0273522|T047|212191006|SNOMEDCT_US|CAUDA EQUINA INJURY WITHOUT BONE INJURY|CAUDA EQUINA INJURY WITHOUT BONY INJURY (DISORDER)
C0273522|T047|212191006|SNOMEDCT_US|CAUDA EQUINA INJURY WITHOUT BONE INJURY |CAUDA EQUINA INJURY WITHOUT BONY INJURY (DISORDER)
C0393841|T047|129617008|SNOMEDCT_US|NEUROPATHY IN LIVER DISEASE|HEPATIC NEUROPATHY (DISORDER)
C0393841|T047|129617008|SNOMEDCT_US|NEUROPATHY IN LIVER DISEASE |HEPATIC NEUROPATHY (DISORDER)
C0393841|T047|129617008|SNOMEDCT_US|HEPATIC NEUROPATHY |HEPATIC NEUROPATHY (DISORDER)
C0393841|T047|129617008|SNOMEDCT_US|HEPATIC NEUROPATHY|HEPATIC NEUROPATHY (DISORDER)
C0160799|T047|23658007|SNOMEDCT_US|LATE EFFECT OF INJURY TO PERIPHERAL NERVE OF SHOULDER GIRDLE AND UPPER LIMB|LATE EFFECT OF INJURY TO PERIPHERAL NERVE OF SHOULDER GIRDLE AND/OR UPPER LIMB
C0160799|T047|23658007|SNOMEDCT_US|SEQUELAE OF INJURY OF NERVE OF UPPER LIMB|LATE EFFECT OF INJURY TO PERIPHERAL NERVE OF SHOULDER GIRDLE AND/OR UPPER LIMB
C0160799|T047|23658007|SNOMEDCT_US|LATE EFFECTS OF INJURY OF PERIPHERAL NERVE OF SHOULDER GIRDLE AND UPPER LIMB |LATE EFFECT OF INJURY TO PERIPHERAL NERVE OF SHOULDER GIRDLE AND/OR UPPER LIMB
C0160799|T047|23658007|SNOMEDCT_US|LATE EFFECTS OF INJURY OF PERIPHERAL NERVE OF SHOULDER GIRDLE AND UPPER LIMB|LATE EFFECT OF INJURY TO PERIPHERAL NERVE OF SHOULDER GIRDLE AND/OR UPPER LIMB
C0160799|T047|23658007|SNOMEDCT_US|LATE EFFECT OF INJURY OF PERIPHERAL NERVE OF SHOULDER GIRDLE AND UPPER LIMB|LATE EFFECT OF INJURY TO PERIPHERAL NERVE OF SHOULDER GIRDLE AND/OR UPPER LIMB
C0160799|T047|23658007|SNOMEDCT_US|LT EFF NERV INJ SHLD/ARM|LATE EFFECT OF INJURY TO PERIPHERAL NERVE OF SHOULDER GIRDLE AND/OR UPPER LIMB
C0160799|T047|23658007|SNOMEDCT_US|LATE EFFECT OF INJURY TO PERIPHERAL NERVE OF SHOULDER GIRDLE AND/OR UPPER LIMB |LATE EFFECT OF INJURY TO PERIPHERAL NERVE OF SHOULDER GIRDLE AND/OR UPPER LIMB
C0160799|T047|23658007|SNOMEDCT_US|LATE EFFECT OF INJURY TO PERIPHERAL NERVE OF SHOULDER GIRDLE AND/OR UPPER LIMB|LATE EFFECT OF INJURY TO PERIPHERAL NERVE OF SHOULDER GIRDLE AND/OR UPPER LIMB
C0270102|T047|206235003|SNOMEDCT_US|BIRTH INJURY TO PERIPHERAL NERVOUS SYSTEM|PERIPHERAL NERVE INJURY DUE TO BIRTH TRAUMA (DISORDER)
C0270102|T047|206235003|SNOMEDCT_US|BIRTH INJURY TO PERIPHERAL NERVOUS SYSTEM, UNSPECIFIED|PERIPHERAL NERVE INJURY DUE TO BIRTH TRAUMA (DISORDER)
C0270102|T047|206235003|SNOMEDCT_US|PERIPHERAL NERVE INJURY DUE TO BIRTH TRAUMA |PERIPHERAL NERVE INJURY DUE TO BIRTH TRAUMA (DISORDER)
C0270102|T047|206235003|SNOMEDCT_US|PERIPHERAL NERVE INJURIES DUE TO BIRTH TRAUMA|PERIPHERAL NERVE INJURY DUE TO BIRTH TRAUMA (DISORDER)
C0270102|T047|206235003|SNOMEDCT_US|PERIPHERAL NERVE INJURY DUE TO BIRTH TRAUMA|PERIPHERAL NERVE INJURY DUE TO BIRTH TRAUMA (DISORDER)
C0270102|T047|206235003|SNOMEDCT_US|PERIPHERAL NERVE INJURY AS BIRTH TRAUMA|PERIPHERAL NERVE INJURY DUE TO BIRTH TRAUMA (DISORDER)
C0270102|T047|206235003|SNOMEDCT_US|PERIPHERAL NERVE INJURY AS BIRTH TRAUMA |PERIPHERAL NERVE INJURY DUE TO BIRTH TRAUMA (DISORDER)
C0270102|T047|206235003|SNOMEDCT_US|PERIPHERAL NERVE INJURY DUE TO BIRTH TRAUMA |PERIPHERAL NERVE INJURY DUE TO BIRTH TRAUMA (DISORDER)
C0270102|T047|206235003|SNOMEDCT_US|BIRTH; INJURY, LACERATION, PERIPHERAL NERVE|PERIPHERAL NERVE INJURY DUE TO BIRTH TRAUMA (DISORDER)
C0270102|T047|206235003|SNOMEDCT_US|BIRTH; INJURY, NERVE, PERIPHERAL|PERIPHERAL NERVE INJURY DUE TO BIRTH TRAUMA (DISORDER)
C0270102|T047|206235003|SNOMEDCT_US|INJURY; BIRTH, LACERATION, PERIPHERAL NERVE|PERIPHERAL NERVE INJURY DUE TO BIRTH TRAUMA (DISORDER)
C0270102|T047|206235003|SNOMEDCT_US|INJURY; BIRTH, NERVE, PERIPHERAL|PERIPHERAL NERVE INJURY DUE TO BIRTH TRAUMA (DISORDER)
C0347066|T047|255128001|SNOMEDCT_US|MALIGNANT INFILTRATION OF PERIPHERAL NERVE|MALIGNANT INFILTRATION OF PERIPHERAL NERVE (DISORDER)
C0347066|T047|255128001|SNOMEDCT_US|NEOPLASM - PNS MALIGNANT INFILTRATION|MALIGNANT INFILTRATION OF PERIPHERAL NERVE (DISORDER)
C0347066|T047|255128001|SNOMEDCT_US|MALIGNANT INFILTRATION OF PERIPHERAL NERVE |MALIGNANT INFILTRATION OF PERIPHERAL NERVE (DISORDER)
C0347066|T047|255128001|SNOMEDCT_US|MALIGNANT INFILTRATION OF PERIPHERAL NERVE |MALIGNANT INFILTRATION OF PERIPHERAL NERVE (DISORDER)
C0270933|T047|21018002|SNOMEDCT_US|INFLAMMATORY NEUROPATHY|INFLAMMATORY NEUROPATHY (DISORDER)
C0270933|T047|21018002|SNOMEDCT_US|INFLAMMATORY NEUROPATHY |INFLAMMATORY NEUROPATHY (DISORDER)
C0270933|T047|21018002|SNOMEDCT_US|INFLAMMATORY NEUROPATHY, NOS|INFLAMMATORY NEUROPATHY (DISORDER)
C0393410|T047|193262003|SNOMEDCT_US|OTHER SPECIFIED DISORDERS OF PERIPHERAL NERVOUS SYSTEM |OTHER SPECIFIED DISORDERS OF PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0393410|T047|193262003|SNOMEDCT_US|OTHER SPECIFIED DISORDERS OF PERIPHERAL NERVOUS SYSTEM|OTHER SPECIFIED DISORDERS OF PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0560607|T047|282742004|SNOMEDCT_US|INTERCOSTAL POST-HERPETIC NEURITIS|INTERCOSTAL POST-HERPETIC NEURITIS (DISORDER)
C0560607|T047|282742004|SNOMEDCT_US|INTERCOSTAL POST-HERPETIC NEURITIS |INTERCOSTAL POST-HERPETIC NEURITIS (DISORDER)
C0582681|T047|304782008|SNOMEDCT_US|LESIONS OF NERVES PLEXUSES AND ROOTS|LESIONS OF NERVES PLEXUSES AND ROOTS (DISORDER)
C0582681|T047|304782008|SNOMEDCT_US|LESIONS OF NERVES PLEXUSES AND ROOTS |LESIONS OF NERVES PLEXUSES AND ROOTS (DISORDER)
C1510429|T047|155085004|SNOMEDCT_US|NEUROPATHIES, ENTRAPMENT|COMPRESSION NEUROPATHY (DISORDER)
C1510429|T047|155085004|SNOMEDCT_US|NEUROPATHY, ENTRAPMENT|COMPRESSION NEUROPATHY (DISORDER)
C1510429|T047|155085004|SNOMEDCT_US|NERVE ENTRAPMENT SYNDROMES|COMPRESSION NEUROPATHY (DISORDER)
C1510429|T047|155085004|SNOMEDCT_US|COMPRESSION NEUROPATHY |COMPRESSION NEUROPATHY (DISORDER)
C1510429|T047|155085004|SNOMEDCT_US|COMPRESSION NEUROPATHY|COMPRESSION NEUROPATHY (DISORDER)
C1510429|T047|155085004|SNOMEDCT_US|ENTRAPMENT NEUROPATHIES|COMPRESSION NEUROPATHY (DISORDER)
C1510429|T047|155085004|SNOMEDCT_US|ENTRAPMENT NEUROPATHY|COMPRESSION NEUROPATHY (DISORDER)
C1510429|T047|155085004|SNOMEDCT_US|NERVE ENTRAPMENT SYNDROME|COMPRESSION NEUROPATHY (DISORDER)
C1510429|T047|155085004|SNOMEDCT_US|TRAPPED NERVE|COMPRESSION NEUROPATHY (DISORDER)
C1510429|T047|155085004|SNOMEDCT_US|PERIPHERAL NERVE ENTRAPMENT SYNDROME |COMPRESSION NEUROPATHY (DISORDER)
C1510429|T047|155085004|SNOMEDCT_US|PERIPHERAL NERVE ENTRAPMENT SYNDROME|COMPRESSION NEUROPATHY (DISORDER)
C1510429|T047|155085004|SNOMEDCT_US|NEUROPATHY; ENTRAPMENT|COMPRESSION NEUROPATHY (DISORDER)
C1510429|T047|155085004|SNOMEDCT_US|ENTRAPMENT SYNDROME, NOS|COMPRESSION NEUROPATHY (DISORDER)
C1510429|T047|155085004|SNOMEDCT_US|ENTRAPMENT NEUROPATHY, NOS|COMPRESSION NEUROPATHY (DISORDER)
C0271684|T047|19378003|SNOMEDCT_US|DIABETIC PSEUDOTABES|DIABETIC PSEUDOTABES (DISORDER)
C0271684|T047|19378003|SNOMEDCT_US|DIABETIC PSEUDOTABES |DIABETIC PSEUDOTABES (DISORDER)
C0564741|T047|286939004|SNOMEDCT_US|OTHER PERIPHERAL NERVE DISEASE|OTHER PERIPHERAL NERVE DISEASE (DISORDER)
C0564741|T047|286939004|SNOMEDCT_US|OTHER PERIPHERAL NERVE DISEASE |OTHER PERIPHERAL NERVE DISEASE (DISORDER)
C3647370|T047||SNOMEDCT_US|NEUROPATHY PERIPHERAL IN ASSOCIATION WITH HEREDITARY ATAXIA 
C3647370|T047||SNOMEDCT_US|NEUROPATHY PERIPHERAL IN ASSOCIATION WITH HEREDITARY ATAXIA
C3662005|T047|609600000|SNOMEDCT_US|NEUROPATHY OF LOWER LIMB|NEUROPATHY OF LOWER LIMB (DISORDER)
C3662005|T047|609600000|SNOMEDCT_US|NEUROPATHY OF LOWER LIMB |NEUROPATHY OF LOWER LIMB (DISORDER)
C1282521|T047|315056009|SNOMEDCT_US|PUDENDAL NERVE NEUROPATHY |PUDENDAL NERVE NEUROPATHY (DISORDER)
C1282521|T047|315056009|SNOMEDCT_US|PUDENDAL NERVE NEUROPATHY|PUDENDAL NERVE NEUROPATHY (DISORDER)
C3662002|T047|609599003|SNOMEDCT_US|NEUROPATHY OF UPPER LIMB |NEUROPATHY OF UPPER LIMB (DISORDER)
C3662002|T047|609599003|SNOMEDCT_US|NEUROPATHY OF UPPER LIMB|NEUROPATHY OF UPPER LIMB (DISORDER)
C3661994|T047|609612001|SNOMEDCT_US|DISORDER OF NERVE ROOT AND/OR PLEXUS |DISORDER OF NERVE ROOT AND/OR PLEXUS (DISORDER)
C3661994|T047|609612001|SNOMEDCT_US|DISORDER OF NERVE ROOT AND/OR PLEXUS|DISORDER OF NERVE ROOT AND/OR PLEXUS (DISORDER)
C0574905|T047|298119007|SNOMEDCT_US|LONG THORACIC NERVE LESION|LONG THORACIC NERVE LESION (DISORDER)
C0574905|T047|298119007|SNOMEDCT_US|LONG THORACIC NERVE LESION |LONG THORACIC NERVE LESION (DISORDER)
C3670522|T047||SNOMEDCT_US|DYSMYELINOGENESIS 
C3670522|T047||SNOMEDCT_US|DYSMYELINOGENESIS
C2931445|T047||SNOMEDCT_US|SACRAL PLEXOPATHY
C1845095|T047||SNOMEDCT_US|DEAFNESS, X-LINKED 5
C1845095|T047||SNOMEDCT_US|DEAFNESS, X-LINKED 5 
C1845095|T047||SNOMEDCT_US|AUDITORY NEUROPATHY, X-LINKED, 1, WITH PERIPHERAL SENSORY NEUROPATHY
C1833831|T047||SNOMEDCT_US|OPTIC ATROPHY, HEARING LOSS, AND PERIPHERAL NEUROPATHY, AUTOSOMAL DOMINANT
C1855885|T047||SNOMEDCT_US|HYPERTROPHIC NEUROPATHY AND CATARACT
C1850383|T047||SNOMEDCT_US|NEUROPATHY, PAINFUL
C1834180|T047||SNOMEDCT_US|NEUROPATHY, WITH PARAPROTEIN IN SERUM, CEREBROSPINAL FLUID AND URINE
C1850022|T047||SNOMEDCT_US|PERIPHERAL NEUROPATHY, ATAXIA, FOCAL NECROTIZING ENCEPHALOPATHY, AND SPONGY DEGENERATION OF BRAIN
C1866770|T047||SNOMEDCT_US|SPINOCEREBELLAR ATAXIA WITH RIGIDITY AND PERIPHERAL NEUROPATHY
C0031315|T047|193115004|SNOMEDCT_US|LIMB, PHANTOM|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|LIMBS, PHANTOM|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PHANTOM LIMB|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PHANTOM LIMBS|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PHANTOM LIMB |PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PHANTOM LIMB SYNDROME WITH PAIN|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PHANTOM LIMB SYNDROME|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PHANTOM LIMB SYNDROME |PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PSEUDOMELIAS|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PHANTOM LIMB SYNDROME NOS|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PHANTOM LIMB [DISEASE/FINDING]|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PSEUDOMELIA|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PHANTOM LIMB SYNDROME WITH PAIN |PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PHANTOM LIMB SYNDROME WITH PAIN |PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PHANTOM LIMB |PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PHANTOM LIMB PAIN|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PLS - PHANTOM LIMB PAIN SYNDROME|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|STUMP HALLUCINATION|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PHANTOM PAIN|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PLS - PHANTOM LIMB SYNDROME|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PHANTOM LIMB SYNDROME |PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|FLS - PHANTOM LIMB SYNDROME|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PAIN; PHANTOM LIMB SYNDROME|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PHANTOM LIMB SYNDROME; PAIN|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PHANTOM LIMB; SYNDROME, WITH PAIN|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|PHANTOM LIMB; SYNDROME|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|SYNDROME; PHANTOM LIMB, WITH PAIN|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C0031315|T047|193115004|SNOMEDCT_US|SYNDROME; PHANTOM LIMB|PHANTOM LIMB SYNDROME WITH PAIN (FINDING)
C3873567|T047|707088000|SNOMEDCT_US|PERIPHERAL NEUROPATHY DUE TO CHEMOTHERAPY|PERIPHERAL NEUROPATHY DUE TO CHEMOTHERAPY (DISORDER)
C3873567|T047|707088000|SNOMEDCT_US|CHEMOTHERAPY-INDUCED PERIPHERAL NEUROPATHY|PERIPHERAL NEUROPATHY DUE TO CHEMOTHERAPY (DISORDER)
C3873567|T047|707088000|SNOMEDCT_US|PERIPHERAL NEUROPATHY DUE TO CHEMOTHERAPY |PERIPHERAL NEUROPATHY DUE TO CHEMOTHERAPY (DISORDER)
C3873567|T047|707088000|SNOMEDCT_US|CIPN - CHEMOTHERAPY-INDUCED PERIPHERAL NEUROPATHY|PERIPHERAL NEUROPATHY DUE TO CHEMOTHERAPY (DISORDER)
C4024907|T047||SNOMEDCT_US|MIXED DEMYELINATING AND AXONAL POLYNEUROPATHY
C0271683|T047|85423005|SNOMEDCT_US|MOTOR POLYNEUROPATHY|MOTOR POLYNEUROPATHY (DISORDER)
C0271683|T047|85423005|SNOMEDCT_US|MOTOR POLYNEUROPATHIES|MOTOR POLYNEUROPATHY (DISORDER)
C0271683|T047|85423005|SNOMEDCT_US|POLYNEUROPATHIES, MOTOR|MOTOR POLYNEUROPATHY (DISORDER)
C0271683|T047|85423005|SNOMEDCT_US|POLYNEUROPATHY, MOTOR|MOTOR POLYNEUROPATHY (DISORDER)
C0271683|T047|85423005|SNOMEDCT_US|MOTOR POLYNEUROPATHY |MOTOR POLYNEUROPATHY (DISORDER)
C1867971|T047||SNOMEDCT_US|ACUTE EPISODES OF NEUROPATHIC SYMPTOMS
C1848695|T047||SNOMEDCT_US|EPISODIC PERIPHERAL NEUROPATHY
C4024974|T047||SNOMEDCT_US|SENSORIMOTOR POLYNEUROPATHY AFFECTING ARMS MORE THAN LEGS
C1112256|T047||SNOMEDCT_US|SENSORIMOTOR PERIPHERAL NEUROPATHY
C1112256|T047||SNOMEDCT_US|PERIPHERAL SENSORIMOTOR NEUROPATHY
C1112256|T047||SNOMEDCT_US|SENSORIMOTOR NEUROPATHY
C1112256|T047||SNOMEDCT_US|MIXED POLYNEUROPATHY
C4024967|T047||SNOMEDCT_US|CONGENITAL PERIPHERAL NEUROPATHY
C4025794|T047||SNOMEDCT_US|CHRONIC SENSORINEURAL POLYNEUROPATHY
C1263857|T047|128208007|SNOMEDCT_US|PERIPHERAL AXONAL NEUROPATHY|PERIPHERAL AXONAL NEUROPATHY (DISORDER)
C1263857|T047|128208007|SNOMEDCT_US|AXONAL PERIPHERAL NEUROPATHY|PERIPHERAL AXONAL NEUROPATHY (DISORDER)
C1263857|T047|128208007|SNOMEDCT_US|PERIPHERAL AXONAL NEUROPATHY |PERIPHERAL AXONAL NEUROPATHY (DISORDER)
C1859178|T047||SNOMEDCT_US|PROGRESSIVE POLYNEUROPATHY
C1859178|T047||SNOMEDCT_US|PROGRESSIVE PERIPHERAL NEUROPATHY
C1859178|T047||SNOMEDCT_US|PERIPHERAL NEUROPATHY, PROGRESSIVE
C4039742|T047|709143008|SNOMEDCT_US|PERIPHERAL NEUROPATHY CAUSED BY TOXIN |PERIPHERAL NEUROPATHY CAUSED BY TOXIN (DISORDER)
C4039742|T047|709143008|SNOMEDCT_US|PERIPHERAL NEUROPATHY CAUSED BY TOXIN|PERIPHERAL NEUROPATHY CAUSED BY TOXIN (DISORDER)
C3495442|T047|247380005|SNOMEDCT_US|PHANTOM PAIN|PHANTOM PAIN (FINDING)
C3495442|T047|247380005|SNOMEDCT_US|PHANTOM PAIN |PHANTOM PAIN (FINDING)
C3495442|T047|247380005|SNOMEDCT_US|PHANTOM LIMB SYNDROME|PHANTOM PAIN (FINDING)
C3495442|T047|247380005|SNOMEDCT_US|PHANTOM PAIN |PHANTOM PAIN (FINDING)
C4039352|T047|709145001|SNOMEDCT_US|PERIPHERAL NEUROPATHY DUE TO INFLAMMATION|PERIPHERAL NEUROPATHY DUE TO INFLAMMATION (DISORDER)
C4039352|T047|709145001|SNOMEDCT_US|PERIPHERAL NEUROPATHY DUE TO INFLAMMATION |PERIPHERAL NEUROPATHY DUE TO INFLAMMATION (DISORDER)
C3276706|T047|709489006|SNOMEDCT_US|SFNP|SFNP - SMALL FIBER NEUROPATHY
C3276706|T047|709489006|SNOMEDCT_US|NEUROPATHY, SMALL FIBER|SFNP - SMALL FIBER NEUROPATHY
C3276706|T047|709489006|SNOMEDCT_US|SMALL FIBRE NEUROPATHY|SFNP - SMALL FIBER NEUROPATHY
C3276706|T047|709489006|SNOMEDCT_US|SMALL FIBER NEUROPATHY|SFNP - SMALL FIBER NEUROPATHY
C3276706|T047|709489006|SNOMEDCT_US|SMALL FIBER NEUROPATHY |SFNP - SMALL FIBER NEUROPATHY
C3276706|T047|709489006|SNOMEDCT_US|SMALL NERVE FIBER NEUROPATHY|SFNP - SMALL FIBER NEUROPATHY
C4040658|T047|710360007|SNOMEDCT_US|PERIPHERAL NEUROPATHY DUE TO METABOLIC DISORDER|PERIPHERAL NEUROPATHY DUE TO METABOLIC DISORDER (DISORDER)
C4040658|T047|710360007|SNOMEDCT_US|PERIPHERAL NEUROPATHY DUE TO METABOLIC DISORDER |PERIPHERAL NEUROPATHY DUE TO METABOLIC DISORDER (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH OR TROCHLEAR NERVE PALSY|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH [TROCHLEAR] NERVE PALSY|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH NERVE PALSY|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH CRANIAL NERVE PALSY|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH NERVE PALSY |FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|IVTH NERVE PARALYSIS|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH NERVE PALSIES|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|PALSIES, FOURTH NERVE|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|PALSY, FOURTH NERVE|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|PALSIES, TROCHLEAR NERVE|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|PALSY, TROCHLEAR NERVE|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|TROCHLEAR NERVE PALSIES|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|TROCHLEAR NERVE DISORDER|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|IVTH CRANIAL NERVE DISORDER|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|TROCHLEAR NERVE DISEASES|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH CRANIAL NERVE DISEASES|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|TROCHLEAR NERVE DISORDERS|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|TROCHLEAR NERVE DISEASES [DISEASE/FINDING]|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|TROCHLEAR NEUROPATHY|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|CRANIAL NERVE IV DISEASES|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|PALSY;IV NERVE|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH CRANIAL NERVE PARESIS |FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|DISORDER OF TROCHLEAR NERVE|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH CRANIAL NERVE DISEASE |FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH CRANIAL NERVE DISEASE|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|SUPERIOR OBLIQUE MUSCLE INNERVATION DISORDER |FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|IVTH NERVE PARESIS|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|SUPERIOR OBLIQUE MUSCLE INNERVATION DISORDER|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|DISORDER OF TROCHLEAR NERVE |FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH CRANIAL NERVE PARESIS|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|DISORDER OF CRANIAL NERVE 4|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|IVTH NERVE DISORDER|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|TROCHLEAR NERVE PALSY|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|SUPERIOR OBLIQUE PALSY|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|TROCHLEAR NERVE PARALYSIS|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|PARESIS OF FOURTH CRANIAL NERVE|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|IVTH NERVE PALSY|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH NERVE PARESIS|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH NERVE PARALYSIS|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH CRANIAL NERVE PARALYSIS|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH CRANIAL NERVE DISORDER|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|TROCHLEAR NERVE WEAKNESS|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|4TH NERVE PALSY|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|IV NERVE PALSY|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH NERVE PALSY |FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|TROCHLEAR NERVE DISEASE|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|DISEASE (OR DISORDER); CRANIAL NERVE, FOURTH|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|DISEASE (OR DISORDER); TROCHLEAR NERVE|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|N.TROCHLEARIS; PARALYSIS|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|PARALYSIS; CRANIAL NERVE, FOURTH|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|PARALYSIS; TROCHLEAR NERVE|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH CRANIAL NERVE DISEASE, NOS|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|FOURTH CRANIAL NERVE DISORDER, NOS|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|TROCHLEAR NERVE DISEASE, NOS|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|TROCHLEAR NERVE DISORDER, NOS|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271375|T047|67883005|SNOMEDCT_US|IV THNERVE PALSY|FOURTH CRANIAL NERVE PARESIS (DISORDER)
C0271353|T047|230531004|SNOMEDCT_US|THIRD CRANIAL NERVE DISORDER|DISORDER OF OCULOMOTOR NERVE (DISORDER)
C0271353|T047|230531004|SNOMEDCT_US|DISORDER OF OCULOMOTOR NERVE|DISORDER OF OCULOMOTOR NERVE (DISORDER)
C0271353|T047|230531004|SNOMEDCT_US|DISORDER OF OCULOMOTOR NERVE |DISORDER OF OCULOMOTOR NERVE (DISORDER)
C0271353|T047|230531004|SNOMEDCT_US|IIIRD NERVE DISORDER|DISORDER OF OCULOMOTOR NERVE (DISORDER)
C0271353|T047|230531004|SNOMEDCT_US|DISORDER OF CRANIAL NERVE 3|DISORDER OF OCULOMOTOR NERVE (DISORDER)
C0271353|T047|230531004|SNOMEDCT_US|OCULOMOTOR NERVE DISORDER|DISORDER OF OCULOMOTOR NERVE (DISORDER)
C0271353|T047|230531004|SNOMEDCT_US|OCULOMOTOR NERVE DISEASE|DISORDER OF OCULOMOTOR NERVE (DISORDER)
C0271353|T047|230531004|SNOMEDCT_US|THIRD CRANIAL NERVE DISEASE |DISORDER OF OCULOMOTOR NERVE (DISORDER)
C0271353|T047|230531004|SNOMEDCT_US|THIRD CRANIAL NERVE DISEASE|DISORDER OF OCULOMOTOR NERVE (DISORDER)
C0271353|T047|230531004|SNOMEDCT_US|CRANIAL NERVE; DISORDER, THIRD (OCULOMOTOR)|DISORDER OF OCULOMOTOR NERVE (DISORDER)
C0271353|T047|230531004|SNOMEDCT_US|DISEASE (OR DISORDER); CRANIAL NERVE, THIRD (OCULOMOTOR)|DISORDER OF OCULOMOTOR NERVE (DISORDER)
C0271353|T047|230531004|SNOMEDCT_US|DISEASE (OR DISORDER); NERVE, OCULOMOTOR|DISORDER OF OCULOMOTOR NERVE (DISORDER)
C0271353|T047|230531004|SNOMEDCT_US|N.OCULOMOTORIUS; DISORDER|DISORDER OF OCULOMOTOR NERVE (DISORDER)
C0271353|T047|230531004|SNOMEDCT_US|OCULOMOTOR NERVE DISEASE, NOS|DISORDER OF OCULOMOTOR NERVE (DISORDER)
C0271353|T047|230531004|SNOMEDCT_US|OCULOMOTOR NERVE DISORDER, NOS|DISORDER OF OCULOMOTOR NERVE (DISORDER)
C0271353|T047|230531004|SNOMEDCT_US|THIRD CRANIAL NERVE DISEASE, NOS|DISORDER OF OCULOMOTOR NERVE (DISORDER)
C0271353|T047|230531004|SNOMEDCT_US|THIRD CRANIAL NERVE DISORDER, NOS|DISORDER OF OCULOMOTOR NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDERS OF PNEUMOGASTRIC (10TH) NERVE|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDERS OF VAGUS NERVE|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|TENTH CRANIAL NERVE DIS|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|PNEUMOGASTRIC NERVE DIS|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|CRANIAL NERVE X DIS|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|VAGUS NERVE DIS|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|VAGUS NERVE DISORDERS|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|VAGUS NERVE DISEASE|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|VAGUS NERVE DISEASES|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDER, PNEUMOGASTRIC NERVE|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDERS, PNEUMOGASTRIC NERVE|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|PNEUMOGASTRIC NERVE DISORDER|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|VAGUS NERVE DISORDER|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|NEUROPATHIES, VAGUS|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|NEUROPATHY, VAGUS|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|VAGUS NEUROPATHIES|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDERS OF PNEUMOGASTRIC [10TH] NERVE|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|TENTH CRANIAL NERVE DISEASES|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|VAGUS NEUROPATHY|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|VAGUS NERVE DISEASES [DISEASE/FINDING]|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|CRANIAL NERVE X DISEASES|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|PNEUMOGASTRIC NERVE DISORDERS|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDER OF VAGUS NERVE |DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDER VAGUS NERVE|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDER OF VAGUS NERVE|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDER OF CRANIAL NERVE 10|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|VAGUS NERVE DISORDER NOS|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDERS OF THE XTH CRANIAL NERVE|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDERS OF THE TENTH NERVE|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|VAGUS NERVE LESION|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDER OF PNEUMOGASTRIC NERVE|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDER OF THE TENTH CRANIAL NERVE|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDER OF VAGUS NERVE |DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|CRANIAL NERVE; DISORDER, TENTH (VAGUS)|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISEASE (OR DISORDER); CRANIAL NERVE, TENTH (VAGUS)|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISEASE (OR DISORDER); NERVE, PNEUMOGASTRIC|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISEASE (OR DISORDER); NERVE, VAGUS|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|N.VAGUS; DISORDER|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDER OF PNEUMOGASTRIC NERVE, NOS|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDER OF THE TENTH CRANIAL NERVE, NOS|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDER OF VAGUS NERVE, NOS|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDER OF PNEUMOGASTRIC NERVE |DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|N.PNEUMOGASTRIC; DISORDER|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDERS OF 10TH NERVE|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDERS OF PNEUMOGASTRIC NERVE|DISORDER OF VAGUS NERVE (DISORDER)
C0152179|T047|73765005|SNOMEDCT_US|DISORDERS OF VAGAL NERVE|DISORDER OF VAGUS NERVE (DISORDER)
C0270923|T047|385006|SNOMEDCT_US|SECONDARY PERIPHERAL NEUROPATHY |SECONDARY PERIPHERAL NEUROPATHY (DISORDER)
C0270923|T047|385006|SNOMEDCT_US|SECONDARY PERIPHERAL NEUROPATHY|SECONDARY PERIPHERAL NEUROPATHY (DISORDER)
C0270923|T047|385006|SNOMEDCT_US|SECONDARY PERIPHERAL NEUROPATHY, NOS|SECONDARY PERIPHERAL NEUROPATHY (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|TRIGEMINAL NERVE DISORDERS|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|DISORDER OF TRIGEMINAL NERVE, UNSPECIFIED|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|DISORDERS OF TRIGEMINAL NERVE|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|CRANIAL NERVE V DIS|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|TRIGEMINAL NERVE DIS|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|FIFTH CRANIAL NERVE DIS|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|TRIGEMINAL DISORDERS|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|TRIGEMINAL NERVE DISEASE|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|TRIGEMINAL NERVE DISEASES|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|TRIGEMINAL NERVE DISORDER|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|NEUROPATHIES, TRIGEMINAL|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|NEUROPATHY, TRIGEMINAL|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|TRIGEMINAL NEUROPATHIES|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|TRIGEMINAL NERVE DIS NOS|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|DISORDERS OF 5TH CRANIAL NERVE|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|TRIGEMINAL NERVE DISEASES [DISEASE/FINDING]|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|CRANIAL NERVE V DISEASES|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|TRIGEMINAL NEUROPATHY|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|FIFTH CRANIAL NERVE DISEASES|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|DISORDER TRIGEMINAL NERVE|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|DISORDER OF TRIGEMINAL NERVE|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|DISORDER OF TRIGEMINAL NERVE |TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|TRIGEMINAL NERVE DISORDER NOS |TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|TRIGEMINAL NERVE DISORDER NOS|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|DISORDER OF TRIGEMINAL NERVE |TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|DISORDER OF CRANIAL NERVE 5|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|TRIGEMINAL NERVE--DISEASES|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|TRIGEMINAL NERVE DISORDER, UNSPECIFIED|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|DISORDERS OF THE VTH CRANIAL NERVE|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|DISORDERS OF THE FIFTH NERVE|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|DISORDER OF THE FIFTH CRANIAL NERVE|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|TRIGEMINAL NERVE DISORDER |TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|DISEASE (OR DISORDER); CRANIAL NERVE, FIFTH|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|DISEASE (OR DISORDER); TRIGEMINAL NERVE|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|DISORDER OF THE FIFTH CRANIAL NERVE, NOS|TRIGEMINAL NERVE DISORDER (DISORDER)
C0152177|T047|64309007|SNOMEDCT_US|TRIGEMINAL NERVE DISORDER, NOS|TRIGEMINAL NERVE DISORDER (DISORDER)
C0031121|T047|25416002|SNOMEDCT_US|PERIPHERAL NEURALGIA|PERIPHERAL NEURALGIA (DISORDER)
C0031121|T047|25416002|SNOMEDCT_US|PERIPHERAL NEURALGIA |PERIPHERAL NEURALGIA (DISORDER)
C4076016|T047|713527009|SNOMEDCT_US|DISORDER OF PERIPHERAL NERVOUS SYSTEM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |DISORDER OF PERIPHERAL NERVOUS SYSTEM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076016|T047|713527009|SNOMEDCT_US|DISORDER OF PERIPHERAL NERVOUS SYSTEM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|DISORDER OF PERIPHERAL NERVOUS SYSTEM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH OR ABDUCENS NERVE PALSY|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH [ABDUCENT] NERVE PALSY|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|LATERAL RECTUS PALSY|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENS NERVE DIS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH CRANIAL NERVE DIS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|VITH CRANIAL NERVE DIS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|CRANIAL NERVE VI DIS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH NERVE PALSY |LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH NERVE PALSY|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH CRANIAL NERVE PALSY|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENS PARALYSIS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|VITH NERVE PARALYSIS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENS NERVE DISEASE|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENS NERVE DISEASES|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENS NERVE PALSIES|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|PALSIES, ABDUCENS NERVE|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|PALSY, ABDUCENS NERVE|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|LATERAL RECTUS PALSIES|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|PALSIES, LATERAL RECTUS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|PALSY, LATERAL RECTUS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|PALSIES, SIXTH NERVE|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|PALSY, SIXTH NERVE|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH NERVE PALSIES|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|PALSY, VI NERVE|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|NERVE PALSIES, VI|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|NERVE PALSY, VI|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|PALSIES, VI NERVE|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|NERVE PALSY, 6TH|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|PALSIES, 6TH NERVE|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|PALSY, 6TH NERVE|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|6TH NERVE PALSIES|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|NERVE PALSIES, 6TH|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENS NERVE PALSY|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|VITH CRANIAL NERVE DISEASES|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|CRANIAL NERVE VI DISEASES|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH CRANIAL NERVE DISORDERS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH CRANIAL NERVE DISEASES|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENS NERVE DISEASES [DISEASE/FINDING]|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|CRANIAL NERVE VI PALSY|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|6TH NERVE PALSY|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|VI NERVE PALSY|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENS NERVE WEAKNESS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH CRANIAL NERVE WEAKNESS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH CRANIAL NERVE DISORDER|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|DISORDER OF ABDUCENT NERVE|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENS (SIXTH) NERVE PALSY|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH CRANIAL NERVE DISEASE|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|DISORDER OF ABDUCENT NERVE |LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|LATERAL RECTUS MUSCLE DENERVATION PARESIS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENS NERVE PARALYSIS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENS NERVE DISORDER|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH CRANIAL NERVE PARALYSIS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|LATERAL RECTUS MUSCLE INNERVATION DISORDER|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|VITH NERVE DISORDER|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|LATERAL RECTUS MUSCLE DENERVATION PARESIS |LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|LATERAL RECTUS MUSCLE INNERVATION DISORDER |LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENS NERVE PARESIS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH CRANIAL NERVE DISEASE |LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH NERVE PALSY |LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|DISORDER OF ABDUCENS NERVE|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|DISORDER OF CRANIAL NERVE 6|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH NERVE PARALYSIS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|VITH NERVE PALSY|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENT NERVE PARALYSIS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENS NERVE DISORDER |LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENS NERVE PALSY |LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENS NERVE WEAKNESS |LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|DISEASE (OR DISORDER); ABDUCENT NERVE|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|DISEASE (OR DISORDER); CRANIAL NERVE, SIXTH|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|PARALYSIS; ABDUCENT NERVE|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|PARALYSIS; CRANIAL NERVE, SIXTH|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENS NERVE DISEASE, NOS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|ABDUCENS NERVE DISORDER, NOS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH CRANIAL NERVE DISEASE, NOS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0271355|T047|4892003|SNOMEDCT_US|SIXTH CRANIAL NERVE DISORDER, NOS|LATERAL RECTUS MUSCLE INNERVATION DISORDER (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|DISORDERS OF GLOSSOPHARYNGEAL NERVE|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|CRANIAL NERVE IX DIS|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|GLOSSOPHARYNGEAL NERVE DIS|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|NINTH CRANIAL NERVE DIS|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|CRANIAL NERVE VIIII DISEASES|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|GLOSSOPHARYNGEAL NERVE DISORDERS|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|GLOSSOPHARYNGEAL NERVE DISEASE|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|GLOSSOPHARYNGEAL NERVE DISEASES|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|CRANIAL NERVE IX DISEASES|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|CRANIAL NERVE IX DISORDERS|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|NINTH CRANIAL NERVE DISEASES|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|GLOSSOPHARYNGEAL NERVE DISEASES [DISEASE/FINDING]|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|DISORDER OF GLOSSOPHARYNGEAL NERVE|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|DISORDER OF GLOSSOPHARYNGEAL NERVE |DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|DISORDER GLOSSOPHARYNGEAL NERVE|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|GLOSSOPHARYNGEAL NERVE DISORDER|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|DISORDER OF CRANIAL NERVE 9|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|GLOSSOPHARYNGEAL NERVE DISORDER NOS|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|DISORDER OF THE NINTH CRANIAL NERVE|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|DISORDER OF IXTH CRANIAL NERVE|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|DISORDER OF NINTH NERVE|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|GLOSSOPHARYNGEAL NERVE LESION|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|DISORDER OF GLOSSOPHARYNGEAL NERVE |DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|CRANIAL NERVE; DISORDER, NINTH (GLOSSOPHARYNGEAL)|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|DISEASE (OR DISORDER); CRANIAL NERVE, NINTH (GLOSSOPHARYNGEAL)|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|DISEASE (OR DISORDER); NERVE, GLOSSOPHARYNGEAL|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|N.GLOSSOPHARYNGEUS; DISORDER|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|IX NERVE DISORDER|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0751941|T047|80962007|SNOMEDCT_US|NINTH NERVE DISORDER|DISORDER OF GLOSSOPHARYNGEAL NERVE (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISEASES, FACIAL NERVE|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL NERVE DISEASE|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL NERVE DISEASES|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL NERVE DISORDERS|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISEASE, FACIAL NERVE|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISORDER OF FACIAL NERVE, UNSPECIFIED|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISORDER OF SEVENTH CRANIAL NERVE|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL NERVE DISORDER|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL NERVE DISORDER |FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL NEUROPATHY|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISORDERS OF THE VIITH CRANIAL NERVE|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISORDERS OF THE SEVENTH NERVE|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISORDER OF FACIAL NERVE|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|SEVENTH CRANIAL NERVE DIS|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|CRANIAL NERVE VII DIS|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL NERVE DIS|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISORDER, FACIAL NERVE|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISORDERS, FACIAL NERVE|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL NEUROPATHIES|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|NEUROPATHIES, FACIAL|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|NEUROPATHY, FACIAL|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL NERVE DIS NOS|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISORDERS OF 7TH CRANIAL NERVE|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|SEVENTH CRANIAL NERVE DISEASES|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|CRANIAL NERVE VII DISORDERS|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL NERVE DISEASES [DISEASE/FINDING]|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|CRANIAL NERVE VII DISEASES|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|LMNL OF VIITH NERVE|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL CRANIAL NERVE DISORDERS|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISORDER OF FACIAL NERVE |FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISORDER FACIAL NERVE|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL NERVE DISORDERS NOS|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL NERVE DISORDER NOS |FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISORDER OF FACIAL NERVE |FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL NERVE DISORDER NOS|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL NEUROPATHY |FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISORDER OF CRANIAL NERVE 7|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL NERVE--DISEASES|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL NERVE DISORDER, UNSPECIFIED|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISEASE (OR DISORDER); CRANIAL NERVE, SEVENTH|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISEASE (OR DISORDER); FACIAL NERVE|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISORDER OF SEVENTH CRANIAL NERVE, NOS|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|FACIAL NERVE DISORDER, NOS|FACIAL NEUROPATHY (DISORDER)
C0015464|T047|230543003|SNOMEDCT_US|DISORDER OF OF SEVENTH CRANIAL NERVE, NOS|FACIAL NEUROPATHY (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISORDERS OF HYPOGLOSSAL (12TH) NERVE|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISORDERS OF HYPOGLOSSAL NERVE|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|HYPOGLOSSAL NERVE DIS|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|CRANIAL NERVE XII DIS|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|TWELFTH CRANIAL NERVE DIS|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|HYPOGLOSSAL NERVE DISORDERS|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|HYPOGLOSSAL NERVE DISEASE|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|HYPOGLOSSAL NERVE DISEASES|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISORDERS OF 12TH CRANIAL NERVE|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|TWELFTH CRANIAL NERVE DISORDER|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|CRANIAL NERVE XII DISEASES|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|CRANIAL NERVE XII DISORDERS|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|HYPOGLOSSAL NERVE DISEASES [DISEASE/FINDING]|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|TWELFTH CRANIAL NERVE DISEASES|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISORDER OF HYPOGLOSSAL NERVE |DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISORDER OF HYPOGLOSSAL NERVE|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISORDER HYPOGLOSSAL NERVE|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|HYPOGLOSSAL NERVE DISORDER|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISORDER OF CRANIAL NERVE 12|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|HYPOGLOSSAL NERVE DISORDER NOS|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISORDERS OF THE XIITH CRANIAL NERVE|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISORDERS OF THE TWELFTH CRANIAL NERVE|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|HYPOGLOSSAL NERVE LESION|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISORDER OF HYPOGLOSSAL NERVE |DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISORDER OF THE TWELFTH CRANIAL NERVE|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|CRANIAL NERVE; DISORDER, TWELFTH (HYPOGLOSSAL)|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISEASE (OR DISORDER); CRANIAL NERVE, TWELFTH (HYPOGLOSSAL)|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISEASE (OR DISORDER); NERVE, HYPOGLOSSAL|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|N.HYPOGLOSSUS; DISORDER|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISORDER OF HYPOGLOSSAL NERVE, NOS|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISORDER OF THE TWELFTH CRANIAL NERVE, NOS|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISORDER OF XII NERVE|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|TWELFTH NERVE DISORDER|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISORDER OF THE XII NERVE|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISORDERS OF HYPOGLOSSAL [12TH] NERVE|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0152181|T047|24777009|SNOMEDCT_US|DISORDERS OF 12TH NERVE|DISORDER OF HYPOGLOSSAL NERVE (DISORDER)
C0266834|T047|20725005|SNOMEDCT_US|FAMILIAL VISCERAL NEUROPATHY|FAMILIAL VISCERAL NEUROPATHY (DISORDER)
C0266834|T047|20725005|SNOMEDCT_US|FAMILIAL VISCERAL NEUROPATHY |FAMILIAL VISCERAL NEUROPATHY (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISORDERS OF ACOUSTIC NERVE|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|VESTIBULOCOCHLEAR NERVE DIS|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|CRANIAL NERVE VIII DIS|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|EIGHTH CRANIAL NERVE DIS|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|AUDITORY NERVE DISORDERS|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|VIIITH CRANIAL NERVE DISORDERS|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|VESTIBULOCOCHLEAR NERVE DISEASE|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|VESTIBULOCOCHLEAR NERVE DISEASES|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|ACOUSTIC NERVE DISORDERS|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|EIGHTH CRANIAL NERVE DISEASES|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|CRANIAL NERVE VIII DISEASES|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|CRANIAL NERVE VIII DISORDERS|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|VESTIBULOCOCHLEAR NERVE DISEASES [DISEASE/FINDING]|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISORDER OF ACOUSTIC NERVE |DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISORDER OF ACOUSTIC NERVE|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|ACOUSTIC NERVE DISORDER NOS|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|ACOUSTIC NERVE DISORDER NOS |DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISORDER OF AUDITORY NERVE|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISORDER OF VESTIBULOCOCHLEAR NERVE|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISORDER OF EIGHTH CRANIAL NERVE|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISORDER OF CRANIAL NERVE 8|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISORDER OF EIGHTH NERVE|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISORDER OF ACOUSTOVESTIBULAR NERVE|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISORDER OF ACOUSTIC NERVE |DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISORDER OF THE VESTIBULOCOCHLEAR NERVE|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|AUDITORY NERVE; DISORDER|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|AUDITORY; NERVE|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|CRANIAL NERVE; DISORDER, EIGHTH (AUDITORY)|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISEASE (OR DISORDER); CRANIAL NERVE, EIGHTH (AUDITORY)|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISEASE (OR DISORDER); NERVE, ACOUSTIC|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISEASE (OR DISORDER); NERVE, AUDITORY|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISORDER; VESTIBULOCOCHLEAR NERVE|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISTURBANCE; VESTIBULOCOCHLEAR NERVE|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|N.VESTIBULOCOCHLEARIS; DISORDER|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISORDER OF ACOUSTIC NERVE, NOS|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISORDER OF EIGHTH NERVE, NOS|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISORDER OF THE VESTIBULOCOCHLEAR NERVE, NOS|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|ACOUSTIC NERVE DISORDER|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|VESTIBULOCOCHLEAR NERVE DISORDER|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0001163|T047|77949003|SNOMEDCT_US|DISORDER OF ACOUSTIC OR EIGHTH NERVE|DISORDER OF ACOUSTIC NERVE (DISORDER)
C0495832|T047||SNOMEDCT_US|INJURY OF PERIPHERAL NERVES OF THORAX
C0495832|T047||SNOMEDCT_US|PERIPHERAL NERVE INJURY OF THORAX 
C0495832|T047||SNOMEDCT_US|PERIPHERAL NERVE INJURY OF THORAX
C0495832|T047||SNOMEDCT_US|PERIPHERAL NERVE INJURY THORAX
C0495832|T047||SNOMEDCT_US|INJURY; NERVE, THORAX, PERIPHERAL
C0677499|T047|443876008|SNOMEDCT_US|RADIAL TUNNEL SYNDROME |SUPINATOR SYNDROME
C0677499|T047|443876008|SNOMEDCT_US|RADIAL TUNNEL SYNDROME|SUPINATOR SYNDROME
C0677499|T047|443876008|SNOMEDCT_US|SUPINATOR SYNDROME|SUPINATOR SYNDROME
C0677499|T047|443876008|SNOMEDCT_US|RADIAL TUNNEL SYNDROME |SUPINATOR SYNDROME
C0677499|T047|443876008|SNOMEDCT_US|RADIAL TUNNEL SYNDROME (SUPINATOR SYNDROME)|SUPINATOR SYNDROME
C0149940|T047|52585001|SNOMEDCT_US|SCIATIC NERVE DIS|SCIATIC NEUROPATHY (DISORDER)
C0149940|T047|52585001|SNOMEDCT_US|NERVE DISEASE, SCIATIC|SCIATIC NEUROPATHY (DISORDER)
C0149940|T047|52585001|SNOMEDCT_US|NERVE DISEASES, SCIATIC|SCIATIC NEUROPATHY (DISORDER)
C0149940|T047|52585001|SNOMEDCT_US|SCIATIC NERVE DISEASE|SCIATIC NEUROPATHY (DISORDER)
C0149940|T047|52585001|SNOMEDCT_US|NEUROPATHIES, SCIATIC|SCIATIC NEUROPATHY (DISORDER)
C0149940|T047|52585001|SNOMEDCT_US|NEUROPATHY, SCIATIC|SCIATIC NEUROPATHY (DISORDER)
C0149940|T047|52585001|SNOMEDCT_US|SCIATIC NEUROPATHIES|SCIATIC NEUROPATHY (DISORDER)
C0149940|T047|52585001|SNOMEDCT_US|SCIATIC NEUROPATHY|SCIATIC NEUROPATHY (DISORDER)
C0149940|T047|52585001|SNOMEDCT_US|SCIATIC NEUROPATHY [DISEASE/FINDING]|SCIATIC NEUROPATHY (DISORDER)
C0149940|T047|52585001|SNOMEDCT_US|SCIATIC NERVE DISEASES|SCIATIC NEUROPATHY (DISORDER)
C0149940|T047|52585001|SNOMEDCT_US|SCIATIC NERVE NEUROPATHY|SCIATIC NEUROPATHY (DISORDER)
C0149940|T047|52585001|SNOMEDCT_US|SCIATIC NERVE--DISEASES|SCIATIC NEUROPATHY (DISORDER)
C0149940|T047|52585001|SNOMEDCT_US|SCIATIC NEUROPATHY |SCIATIC NEUROPATHY (DISORDER)
C0149940|T047|52585001|SNOMEDCT_US|DISEASE (OR DISORDER); NERVE, SCIATIC|SCIATIC NEUROPATHY (DISORDER)
C0149940|T047|52585001|SNOMEDCT_US|N.ISCHIADICUS; NEUROPATHIC|SCIATIC NEUROPATHY (DISORDER)
C0149940|T047|52585001|SNOMEDCT_US|NEUROPATHY; SCIATIC NERVE|SCIATIC NEUROPATHY (DISORDER)
C0027881|T047||SNOMEDCT_US|NEURONITIS
C0393804|T047|193197008|SNOMEDCT_US|POLYNEUROPATHY IN DISEASE NOS |POLYNEUROPATHY IN DISEASE NOS (DISORDER)
C0393804|T047|193197008|SNOMEDCT_US|POLYNEUROPATHY IN DISEASE NOS|POLYNEUROPATHY IN DISEASE NOS (DISORDER)
C0477401|T047|194528005|SNOMEDCT_US|OTHER DISORDERS OF PERIPHERAL NERVOUS SYSTEM|[X]OTHER DISORDERS OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0477401|T047|194528005|SNOMEDCT_US|[X]OTHER DISORDERS OF THE PERIPHERAL NERVOUS SYSTEM|[X]OTHER DISORDERS OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0477401|T047|194528005|SNOMEDCT_US|[X]OTHER DISORDERS OF THE PERIPHERAL NERVOUS SYSTEM |[X]OTHER DISORDERS OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0392555|T047|18708008|SNOMEDCT_US|HYPERTROPHIC INTERSTITIAL NEUROPATHY|HYPERTROPHIC INTERSTITIAL NEUROPATHY (DISORDER)
C0392555|T047|18708008|SNOMEDCT_US|HYPERTROPHIC INTERSTITIAL NEUROPATHY |HYPERTROPHIC INTERSTITIAL NEUROPATHY (DISORDER)
C0263899|T047|69071001|SNOMEDCT_US|RADICULAR SYNDROME OF LOWER LIMBS|RADICULAR SYNDROME OF LOWER LIMBS (DISORDER)
C0263899|T047|69071001|SNOMEDCT_US|RADICULAR SYNDROME OF LOWER LIMBS |RADICULAR SYNDROME OF LOWER LIMBS (DISORDER)
C0271348|T047|75834006|SNOMEDCT_US|STRACHAN'S SYNDROME|STRACHAN'S SYNDROME (DISORDER)
C0271348|T047|75834006|SNOMEDCT_US|STRACHAN'S SYNDROME |STRACHAN'S SYNDROME (DISORDER)
C0271348|T047|75834006|SNOMEDCT_US|STRACHAN SYNDROME|STRACHAN'S SYNDROME (DISORDER)
C0271348|T047|75834006|SNOMEDCT_US|AMBLYOPIA, NEUROPATHY, OROGENITAL DERMATITIS SYNDROME|STRACHAN'S SYNDROME (DISORDER)
C0271348|T047|75834006|SNOMEDCT_US|HOWES-PALLISTER-LANDOR SYNDROME|STRACHAN'S SYNDROME (DISORDER)
C0271348|T047|75834006|SNOMEDCT_US|STRACHAN'S SYNDROME |STRACHAN'S SYNDROME (DISORDER)
C0266513|T047|204080008|SNOMEDCT_US|DEFECTIVE DEVELOPMENT OF CAUDA EQUINA|DEFECTIVE DEVELOPMENT OF THE CAUDA EQUINA (DISORDER)
C0266513|T047|204080008|SNOMEDCT_US|DEFECTIVE DEVELOPMENT OF CAUDA EQUINA |DEFECTIVE DEVELOPMENT OF THE CAUDA EQUINA (DISORDER)
C0266513|T047|204080008|SNOMEDCT_US|DEFECTIVE DEVELOPMENT OF THE CAUDA EQUINA|DEFECTIVE DEVELOPMENT OF THE CAUDA EQUINA (DISORDER)
C0266513|T047|204080008|SNOMEDCT_US|DEFECTIVE DEVELOPMENT OF THE CAUDA EQUINA |DEFECTIVE DEVELOPMENT OF THE CAUDA EQUINA (DISORDER)
C0266513|T047|204080008|SNOMEDCT_US|DEVELOPMENT; DEFECTIVE, CONGENITAL, CAUDA EQUINA|DEFECTIVE DEVELOPMENT OF THE CAUDA EQUINA (DISORDER)
C0394022|T047|230803002|SNOMEDCT_US|DISORDER OF NERVE REPAIR|DISORDER OF NERVE REPAIR (DISORDER)
C0394022|T047|230803002|SNOMEDCT_US|DISORDER OF NERVE REPAIR |DISORDER OF NERVE REPAIR (DISORDER)
C0393866|T047|230613008|SNOMEDCT_US|INJECTION NEUROPATHY|INJECTION NEUROPATHY (DISORDER)
C0393866|T047|230613008|SNOMEDCT_US|INJECTION NEUROPATHY |INJECTION NEUROPATHY (DISORDER)
C0555208|T047|253192007|SNOMEDCT_US|FIBROLIPOMA OF FILUM TERMINALE|FIBROLIPOMA OF FILUM TERMINALE (DISORDER)
C0555208|T047|253192007|SNOMEDCT_US|FIBROLIPOMA OF FILUM TERMINALE |FIBROLIPOMA OF FILUM TERMINALE (DISORDER)
C0266516|T047|22133005|SNOMEDCT_US|CONGENITAL MALFORMATIONS ANOMALY OF PERIPHERAL NERVOUS SYSTEM|CONGENITAL ANOMALY OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0266516|T047|22133005|SNOMEDCT_US|CONGENITAL ANOMALY OF PERIPHERAL NERVOUS SYSTEM|CONGENITAL ANOMALY OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0266516|T047|22133005|SNOMEDCT_US|CONGENITAL ANOMALY OF PERIPHERAL NERVOUS SYSTEM |CONGENITAL ANOMALY OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0266516|T047|22133005|SNOMEDCT_US|CONGENITAL PERIPHERAL NERVOUS SYSTEM ANOMALY NOS|CONGENITAL ANOMALY OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0266516|T047|22133005|SNOMEDCT_US|CONGENITAL ANOMALY OF THE PERIPHERAL NERVOUS SYSTEM |CONGENITAL ANOMALY OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0266516|T047|22133005|SNOMEDCT_US|CONGENITAL ANOMALY OF THE PERIPHERAL NERVOUS SYSTEM|CONGENITAL ANOMALY OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C0266516|T047|22133005|SNOMEDCT_US|CONGENITAL ANOMALY OF THE PERIPHERAL NERVOUS SYSTEM, NOS|CONGENITAL ANOMALY OF THE PERIPHERAL NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|ANS DISEASE|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC NERVOUS SYSTEM DISEASES|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|DISORDERS OF THE AUTONOMIC NERVOUS SYSTEM|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC DISEASE|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|DISORDER OF AUTONOMIC NERVOUS SYSTEM, UNSPECIFIED|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|DISORDERS OF AUTONOMIC NERVOUS SYSTEM|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC DISORDER|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC DYSFUNCTION|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|DIS AUTONOMIC NERVOUS SYSTEM|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC NERVOUS SYSTEM DIS|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|ANS DIS|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|NERVOUS SYSTEM DIS AUTONOMIC|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|CENTRAL AUTONOMIC NERVOUS SYSTEM DIS|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC DIS|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC NERVOUS SYSTEM DISORDER |DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC NERVOUS SYSTEM DISORDER|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|ANS DISORDER|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC NERVOUS SYSTEM DISORDERS|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC NERVE DIS NEC|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|DISORDER OF THE AUTONOMIC NERVOUS SYSTEM, UNSPECIFIED|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC CENTRAL NERVOUS SYSTEM DISEASES|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC NERVOUS SYSTEM DISEASES [DISEASE/FINDING]|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|ANS DISEASES|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC DISEASES|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|NERVOUS SYSTEM DISEASES, AUTONOMIC|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|CENTRAL AUTONOMIC NERVOUS SYSTEM DISEASES|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|ANS (AUTONOMIC NERVOUS SYSTEM) DISEASES|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC CNS DIS|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC NERVOUS SYSTEM DISORDER NOS |DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC NERVOUS SYSTEM DISORDER NOS|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC NERVOUS SYSTEM--DISEASES|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|UNSPECIFIED DISORDER OF AUTONOMIC NERVOUS SYSTEM|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|DISORDER OF AUTONOMIC NERVOUS SYSTEM |DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|DISORDER OF AUTONOMIC NERVOUS SYSTEM|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|DISORDER OF VEGETATIVE SYSTEM|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|AUTONOMIC; NERVOUS SYSTEM, DISORDER|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|DISEASE (OR DISORDER); AUTONOMIC NERVOUS SYSTEM|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|DISEASE (OR DISORDER); NERVOUS SYSTEM, AUTONOMIC|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|DISEASE (OR DISORDER); NERVOUS SYSTEM, VEGETATIVE|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|NERVOUS SYSTEM; DISORDER, AUTONOMIC|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|DISORDER OF AUTONOMIC NERVOUS SYSTEM, NOS|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1145628|T047|15241006|SNOMEDCT_US|DISORDER OF VEGETATIVE SYSTEM, NOS|DISORDER OF AUTONOMIC NERVOUS SYSTEM (DISORDER)
C1278821|T047|180234006|SNOMEDCT_US|INFECTIOUS DISORDER OF THE PERIPHERAL NERVOUS SYSTEM|INFECTIOUS PERIPHERAL NEUROPATHY
C1278821|T047|180234006|SNOMEDCT_US|INFECTIOUS DISORDER OF THE PERIPHERAL NERVOUS SYSTEM |INFECTIOUS PERIPHERAL NEUROPATHY
C1278821|T047|180234006|SNOMEDCT_US|PERIPHERAL NERVE INFECTION|INFECTIOUS PERIPHERAL NEUROPATHY
C1278821|T047|180234006|SNOMEDCT_US|INFECTIOUS PERIPHERAL NEUROPATHY|INFECTIOUS PERIPHERAL NEUROPATHY
C1278821|T047|180234006|SNOMEDCT_US|INFECTIOUS DISORDER OF THE PERIPHERAL NERVOUS SYSTEM [AMBIGUOUS]|INFECTIOUS PERIPHERAL NEUROPATHY
C1278821|T047|180234006|SNOMEDCT_US|PERIPHERAL NERVOUS SYSTEM INFECTIOUS DISORDER|INFECTIOUS PERIPHERAL NEUROPATHY
C0270891|T047|2231001|SNOMEDCT_US|ELECTROPHYS: NERVE PLEXUS DISORDER|NERVE PLEXUS DISORDER (DISORDER)
C0270891|T047|2231001|SNOMEDCT_US|NERVE PLEXUS DISORDER |NERVE PLEXUS DISORDER (DISORDER)
C0270891|T047|2231001|SNOMEDCT_US|NERVE PLEXUS DISORDER|NERVE PLEXUS DISORDER (DISORDER)
C0270891|T047|2231001|SNOMEDCT_US|NERVE PLEXUS DISORDER, NOS|NERVE PLEXUS DISORDER (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|DYSTROPHIES, REFLEX SYMPATHETIC|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|DYSTROPHY, REFLEX SYMPATHETIC|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|REFLEX SYMPATHETIC DYSTROPHIES|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|REFLEX SYMPATHETIC DYSTROPHY|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SHOULDER HAND SYNDROME|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SUDECK'S ATROPHY|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SYMPATHETIC DYSTROPHIES, REFLEX|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SYMPATHETIC DYSTROPHY, REFLEX|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SYNDROME, SHOULDER-HAND|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SHOULDER-HAND SYNDROMES|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SYNDROMES, SHOULDER-HAND|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|CRPS TYPE I|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|REFLEX SYMPATHETIC DYSTROPHY OF UPPER EXTREMITY|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SUDECK'S ATROPHY |SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SHOULDER-HAND SYNDROME |SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SHOULDER-HAND SYNDROME|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|COMPLEX REGIONAL PAIN SYNDROME TYPE I OF THE UPPER LIMB|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|ATROPHY, SUDEK|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|ATROPHY, SUDEK'S|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SUDEKS ATROPHY|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|I, CPRS TYPE|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|TYPE I, CPRS|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|REFLEX DYSTROPHIA, SYMPATHETIC|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SYMPATHETIC REFLEX DYSTROPHIAS|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|UNSP RFLX SYMPTH DYSTRPH|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|RFLX SYM DYSTRPH UP LIMB|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SUDEK'S ATROPHY|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|CPRS TYPE I|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|PAIN SYNDROME TYPE I, REGIONAL, COMPLEX|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|COMPLEX REGIONAL PAIN SYNDROME, TYPE I|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|RSD (REFLEX SYMPATHETIC DYSTROPHY)|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SYNDROME, REFLEX SYMPATHETIC DYSTROPHY|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SYMPATHETIC REFLEX DYSTROPHIA|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|TYPE I COMPLEX REGIONAL PAIN SYNDROME|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|REFLEX SYMPATHETIC DYSTROPHY [DISEASE/FINDING]|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|PAIN SYNDROME TYPE I, COMPLEX REGIONAL|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|REFLEX SYMPATHETIC DYSTROPHY SYNDROME|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SUDEK ATROPHY|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|DYSTROPHY;REFLEX SYMPATHETIC|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|ATROPHIES, SUDEK'S|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|CPRS TYPE IS|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|IS, CPRS TYPE|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|RSDS (REFLEX SYMPATHETIC DYSTROPHY)|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SUDEK'S ATROPHIES|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|TYPE IS, CPRS|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|ALGODYSTROPHY|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SUDECK'S ATROPHY |SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|REFLEX SYMPATHETIC DYSTROPHY |SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|REFLEX SYMPATHETIC DYSTROPHY (& SUDEK'S ATROPHY) |SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|CRPS - COMPLEX REGIONAL PAIN SYNDROME TYPE I|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|REFLEX SYMPATHETIC DYSTROPHY (& SUDEK'S ATROPHY)|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SUDEK'S ATROPHY |SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SHOULDER-HAND SYNDROME |SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|RSD - REFLEX SYMPATHETIC DYSTROPHY|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|COMPLEX REGIONAL PAIN SYNDROME TYPE I|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|ALGONEURODYSTROPHY|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|COMPLEX REGIONAL PAIN SYNDROME TYPE I OF UPPER LIMB |SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|COMPLEX REGIONAL PAIN SYNDROME TYPE I |SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|COMPLEX REGIONAL PAIN SYNDROME TYPE I OF UPPER LIMB|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|REFLEX SYMPATHETIC DYSTROPHY OF THE UPPER LIMB|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|REFLEX SYMPATHETIC DYSTROPHY, UNSPECIFIED|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|REFLEX NEUROVASCULAR DYSTROPHY|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|CRPS I|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|RND|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|RSDS|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|COMPLEX REGIONAL PAIN SYNDROME I|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|STEINBROCKER'S SYNDROME|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|ALGODYSTROPHY |SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|REFLEX SYMPATHETIC DYSTROPHY OF UPPER EXTREMITY |SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|ATROPHY; SUDECK|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SUDECK; ATROPHY|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SUDECK|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|HAND-SHOULDER; SYNDROME|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SHOULDER-HAND; SYNDROME|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SYNDROME; HAND-SHOULDER|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|SYNDROME; SHOULDER-HAND|SUDECK'S ATROPHY (DISORDER)
C0034931|T047|156849009|SNOMEDCT_US|REFLEX SYMPATHETIC DYSTROPHY [AMBIGUOUS]|SUDECK'S ATROPHY (DISORDER)
C0494493|T047||SNOMEDCT_US|IDIOPATHIC PROGRESSIVE NEUROPATHY
C0494493|T047||SNOMEDCT_US|IDIOPATHIC PERIPHERAL NEUROPATHY PROGRESSIVE
C0494493|T047||SNOMEDCT_US|IDIOPATHIC PROGRESSIVE NEUROPATHY 
C0494493|T047||SNOMEDCT_US|IDIOPATHIC; NEUROPATHIC, PROGRESSIVE
C0494493|T047||SNOMEDCT_US|NEUROPATHY; IDIOPATHIC, PROGRESSIVE
C0086957|T047|54995001|SNOMEDCT_US|SCALENUS ANTICUS SYNDROME|CERVICAL RIB SYNDROME (DISORDER)
C0086957|T047|54995001|SNOMEDCT_US|SYNDROME, SCALENUS ANTICUS|CERVICAL RIB SYNDROME (DISORDER)
C0086957|T047|54995001|SNOMEDCT_US|SCALENUS ANTICUS SYNDROME |CERVICAL RIB SYNDROME (DISORDER)
C0086957|T047|54995001|SNOMEDCT_US|CERVICAL RIB SYNDROME|CERVICAL RIB SYNDROME (DISORDER)
C0086957|T047|54995001|SNOMEDCT_US|CERVICAL RIB SYNDROME |CERVICAL RIB SYNDROME (DISORDER)
C0086957|T047|54995001|SNOMEDCT_US|SCALENUS ANTICUS SYNDROME |CERVICAL RIB SYNDROME (DISORDER)
C0086957|T047|54995001|SNOMEDCT_US|SCALENUS ANTICUS; SYNDROME|CERVICAL RIB SYNDROME (DISORDER)
C0086957|T047|54995001|SNOMEDCT_US|SYNDROME; SCALENUS ANTICUS|CERVICAL RIB SYNDROME (DISORDER)
C0086957|T047|54995001|SNOMEDCT_US|NAFFZIGER'S SYNDROME|CERVICAL RIB SYNDROME (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|POSTERIOR TIBIAL NERVE DIS|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|TIBIAL NERVE DIS|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|NERVE DISEASE, TIBIAL|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|NERVE DISEASES, TIBIAL|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|TIBIAL NERVE DISEASE|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|INTERNAL POPLITEAL NEUROPATHIES|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|NEUROPATHIES, INTERNAL POPLITEAL|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|NEUROPATHY, INTERNAL POPLITEAL|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|POPLITEAL NEUROPATHIES, INTERNAL|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|POPLITEAL NEUROPATHY, INTERNAL|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|MEDIAL POPLITEAL NEUROPATHIES|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|NEUROPATHIES, MEDIAL POPLITEAL|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|NEUROPATHY, MEDIAL POPLITEAL|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|POPLITEAL NEUROPATHIES, MEDIAL|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|POPLITEAL NEUROPATHY, MEDIAL|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|NEUROPATHIES, POSTERIOR TIBIAL|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|NEUROPATHY, POSTERIOR TIBIAL|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|POSTERIOR TIBIAL NEUROPATHIES|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|TIBIAL NEUROPATHIES, POSTERIOR|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|TIBIAL NEUROPATHY, POSTERIOR|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|NEUROPATHIES, TIBIAL|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|NEUROPATHY, TIBIAL|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|TIBIAL NEUROPATHIES|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|TIBIAL NEUROPATHY|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|TIBIAL NERVE DISEASES|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|TIBIAL NEUROPATHY [DISEASE/FINDING]|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|INTERNAL POPLITEAL NEUROPATHY|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|POSTERIOR TIBIAL NERVE DISEASES|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|POSTERIOR TIBIAL NEUROPATHY|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|MEDIAL POPLITEAL NEUROPATHY|TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|TIBIAL NEUROPATHY |TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|POSTERIOR TIBIAL NEUROPATHY |TIBIAL NEUROPATHY (DISORDER)
C0751932|T047|399076001|SNOMEDCT_US|TIBIAL NEUROPATHY  [AMBIGUOUS]|TIBIAL NEUROPATHY (DISORDER)
C1275816|T047|399088004|SNOMEDCT_US|COMMON PERONEAL NERVE PARALYSIS|COMMON PERONEAL NERVE PARALYSIS (DISORDER)
C1275816|T047|399088004|SNOMEDCT_US|COMMON PERONEAL NERVE PARALYSIS |COMMON PERONEAL NERVE PARALYSIS (DISORDER)
C0205930|T047|7359008|SNOMEDCT_US|ALGONEURODYSTROPHY|ALGONEURODYSTROPHY (DISORDER)
C0205930|T047|7359008|SNOMEDCT_US|ALGONEURODYSTROPHY, UNSPECIFIED SITE|ALGONEURODYSTROPHY (DISORDER)
C0205930|T047|7359008|SNOMEDCT_US|ALGONEURODYSTROPHY NOS|ALGONEURODYSTROPHY (DISORDER)
C0205930|T047|7359008|SNOMEDCT_US|ALGONEURODYSTROPHY NOS |ALGONEURODYSTROPHY (DISORDER)
C0205930|T047|7359008|SNOMEDCT_US|ALGONEURODYSTROPHY |ALGONEURODYSTROPHY (DISORDER)
C0434564|T047|209086000|SNOMEDCT_US|CLOSED DISLOCATION OF LUMBAR VERTEBRA WITH CAUDA EQUINA LESION |CLOSED SPINAL DISLOCATION WITH CAUDA EQUINA LESION (DISORDER)
C0434564|T047|209086000|SNOMEDCT_US|CLOSED DISLOCATION OF LUMBAR VERTEBRA WITH CAUDA EQUINA LESION|CLOSED SPINAL DISLOCATION WITH CAUDA EQUINA LESION (DISORDER)
C0434564|T047|209086000|SNOMEDCT_US|DISLOCATION VERTEBRA LUMBAR CLOSED WITH CAUDA EQUINA LESION|CLOSED SPINAL DISLOCATION WITH CAUDA EQUINA LESION (DISORDER)
C0434564|T047|209086000|SNOMEDCT_US|CLOSED SPINAL DISLOCATION WITH CAUDA EQUINA LESION|CLOSED SPINAL DISLOCATION WITH CAUDA EQUINA LESION (DISORDER)
C0434564|T047|209086000|SNOMEDCT_US|CLOSED SPINAL DISLOCATION WITH CAUDA EQUINA LESION |CLOSED SPINAL DISLOCATION WITH CAUDA EQUINA LESION (DISORDER)
C0434571|T047|209102002|SNOMEDCT_US|OPEN DISLOCATION OF LUMBAR VERTEBRA WITH CAUDA EQUINA LESION|OPEN SPINAL DISLOCATION WITH CAUDA EQUINA LESION (DISORDER)
C0434571|T047|209102002|SNOMEDCT_US|DISLOCATION VERTEBRA OPEN WITH CAUDA EQUINA LESION|OPEN SPINAL DISLOCATION WITH CAUDA EQUINA LESION (DISORDER)
C0434571|T047|209102002|SNOMEDCT_US|OPEN DISLOCATION OF LUMBAR VERTEBRA WITH CAUDA EQUINA LESION |OPEN SPINAL DISLOCATION WITH CAUDA EQUINA LESION (DISORDER)
C0434571|T047|209102002|SNOMEDCT_US|DISLOCATION VERTEBRA LUMBAR OPEN WITH CAUDA EQUINA LESION|OPEN SPINAL DISLOCATION WITH CAUDA EQUINA LESION (DISORDER)
C0434571|T047|209102002|SNOMEDCT_US|OPEN DISLOCATION OF VERTEBRA WITH CAUDA EQUINA LESION|OPEN SPINAL DISLOCATION WITH CAUDA EQUINA LESION (DISORDER)
C0434571|T047|209102002|SNOMEDCT_US|OPEN SPINAL DISLOCATION WITH CAUDA EQUINA LESION|OPEN SPINAL DISLOCATION WITH CAUDA EQUINA LESION (DISORDER)
C0434571|T047|209102002|SNOMEDCT_US|OPEN SPINAL DISLOCATION WITH CAUDA EQUINA LESION |OPEN SPINAL DISLOCATION WITH CAUDA EQUINA LESION (DISORDER)
C0270907|T047|4724003|SNOMEDCT_US|ACUTE RADIAL NERVE PALSY|ACUTE RADIAL NERVE PALSY (DISORDER)
C0270907|T047|4724003|SNOMEDCT_US|ACUTE RADIAL NERVE PALSY |ACUTE RADIAL NERVE PALSY (DISORDER)
C0751922|T047|397828008|SNOMEDCT_US|MEDIAN NEUROPATHY |MEDIAN NEUROPATHY (FINDING)
C0751922|T047|397828008|SNOMEDCT_US|MEDIAN NERVE DIS|MEDIAN NEUROPATHY (FINDING)
C0751922|T047|397828008|SNOMEDCT_US|NERVE PALSY MEDIAN|MEDIAN NEUROPATHY (FINDING)
C0751922|T047|397828008|SNOMEDCT_US|MEDIAN NERVE PALSY|MEDIAN NEUROPATHY (FINDING)
C0751922|T047|397828008|SNOMEDCT_US|MEDIAN NERVE PALSY |MEDIAN NEUROPATHY (FINDING)
C0751922|T047|397828008|SNOMEDCT_US|MEDIAN NERVE DISEASE|MEDIAN NEUROPATHY (FINDING)
C0751922|T047|397828008|SNOMEDCT_US|NERVE DISEASE, MEDIAN|MEDIAN NEUROPATHY (FINDING)
C0751922|T047|397828008|SNOMEDCT_US|NERVE DISEASES, MEDIAN|MEDIAN NEUROPATHY (FINDING)
C0751922|T047|397828008|SNOMEDCT_US|MEDIAN NEUROPATHIES|MEDIAN NEUROPATHY (FINDING)
C0751922|T047|397828008|SNOMEDCT_US|MEDIAN NEUROPATHY|MEDIAN NEUROPATHY (FINDING)
C0751922|T047|397828008|SNOMEDCT_US|NEUROPATHIES, MEDIAN|MEDIAN NEUROPATHY (FINDING)
C0751922|T047|397828008|SNOMEDCT_US|NEUROPATHY, MEDIAN|MEDIAN NEUROPATHY (FINDING)
C0751922|T047|397828008|SNOMEDCT_US|MEDIAN NERVE DISEASES|MEDIAN NEUROPATHY (FINDING)
C0751922|T047|397828008|SNOMEDCT_US|MEDIAN NEUROPATHY [DISEASE/FINDING]|MEDIAN NEUROPATHY (FINDING)
C0751922|T047|397828008|SNOMEDCT_US|MEDIAN NEUROPATHY |MEDIAN NEUROPATHY (FINDING)
C0751922|T047|397828008|SNOMEDCT_US|DISEASE (OR DISORDER); MEDIAN NERVE|MEDIAN NEUROPATHY (FINDING)
C0740447|T047|424736006|SNOMEDCT_US|DIABETIC PERIPHERAL NEUROPATHY |DIABETIC PERIPHERAL NEUROPATHY (DISORDER)
C0740447|T047|424736006|SNOMEDCT_US|DIABETIC PERIPHERAL NEUROPATHY|DIABETIC PERIPHERAL NEUROPATHY (DISORDER)
C0740447|T047|424736006|SNOMEDCT_US|DIABETIC PERIPHERAL NEUROPATHY |DIABETIC PERIPHERAL NEUROPATHY (DISORDER)
C0553761|T047|193129003|SNOMEDCT_US|MEDIAN NERVE COMPRESSION IN FOREARM|MEDIAN NERVE COMPRESSION IN FOREARM (DISORDER)
C0553761|T047|193129003|SNOMEDCT_US|MEDIAN NERVE COMPRESSION IN FOREARM |MEDIAN NERVE COMPRESSION IN FOREARM (DISORDER)
C1384669|T047|399088004|SNOMEDCT_US|LATERAL POPLITEAL NERVE PALSY |COMMON PERONEAL NERVE PALSY
C1384669|T047|399088004|SNOMEDCT_US|NERVE PALSY LATERAL POPLITEAL|COMMON PERONEAL NERVE PALSY
C1384669|T047|399088004|SNOMEDCT_US|NERVE PALSY COMMON PERONEAL|COMMON PERONEAL NERVE PALSY
C1384669|T047|399088004|SNOMEDCT_US|COMMON PERONEAL NERVE PALSY|COMMON PERONEAL NERVE PALSY
C1384669|T047|399088004|SNOMEDCT_US|LATERAL POPLITEAL NERVE PALSY|COMMON PERONEAL NERVE PALSY
C1384669|T047|399088004|SNOMEDCT_US|COMMON PERONEAL NERVE PALSY |COMMON PERONEAL NERVE PALSY
C1335029|T047||SNOMEDCT_US|NON-NEOPLASTIC PERIPHERAL NERVOUS SYSTEM DISEASE
C1335029|T047||SNOMEDCT_US|NON-NEOPLASTIC PERIPHERAL NERVOUS SYSTEM DISORDER
C0026849|T047|193260006|SNOMEDCT_US|MUSCULAR DYSTROPHIES AND OTHER MYOPATHIES|OTHER MYOPATHIES AND MUSCULAR DYSTROPHIES (DISORDER)
C0026849|T047|193260006|SNOMEDCT_US|OTHER MUSCULAR DYSTROPHIES AND MYOPATHIES|OTHER MYOPATHIES AND MUSCULAR DYSTROPHIES (DISORDER)
C0026849|T047|193260006|SNOMEDCT_US|MUSCULAR DYSTROPHIES AND OTHER MYOPATHIES, UNSPECIFIED|OTHER MYOPATHIES AND MUSCULAR DYSTROPHIES (DISORDER)
C0026849|T047|193260006|SNOMEDCT_US|MUSCULAR DYSTROPHY/MYOPATHIES|OTHER MYOPATHIES AND MUSCULAR DYSTROPHIES (DISORDER)
C0026849|T047|193260006|SNOMEDCT_US|OTHER MYOPATHIES AND MUSCULAR DYSTROPHIES|OTHER MYOPATHIES AND MUSCULAR DYSTROPHIES (DISORDER)
C0026849|T047|193260006|SNOMEDCT_US|OTHER MYOPATHIES AND MUSCULAR DYSTROPHIES |OTHER MYOPATHIES AND MUSCULAR DYSTROPHIES (DISORDER)
C0026849|T047|193260006|SNOMEDCT_US|MUSCULAR DYSTROPHIES AND OTHER MYOPATHIES |OTHER MYOPATHIES AND MUSCULAR DYSTROPHIES (DISORDER)
C0154730|T047|193098000|SNOMEDCT_US|DISORDERS OF OTHER CRANIAL NERVES|OTHER CRANIAL NERVE DISORDERS (DISORDER)
C0154730|T047|193098000|SNOMEDCT_US|OTHER CRANIAL NERVE DISORDERS|OTHER CRANIAL NERVE DISORDERS (DISORDER)
C0154730|T047|193098000|SNOMEDCT_US|OTHER CRANIAL NERVE DISORDERS |OTHER CRANIAL NERVE DISORDERS (DISORDER)
C0154747|T047|193154003|SNOMEDCT_US|MONONEURITIS OF LOWER LIMB |UNSPECIFIED MONONEURITIS LOWER LIMB (DISORDER)
C0154747|T047|193154003|SNOMEDCT_US|MONONEURITIS LOWER LIMB|UNSPECIFIED MONONEURITIS LOWER LIMB (DISORDER)
C0154747|T047|193154003|SNOMEDCT_US|MONONEURITIS OF LOWER LIMB|UNSPECIFIED MONONEURITIS LOWER LIMB (DISORDER)
C0154747|T047|193154003|SNOMEDCT_US|MONONEURITIS OF A LOWER LIMB|UNSPECIFIED MONONEURITIS LOWER LIMB (DISORDER)
C0154747|T047|193154003|SNOMEDCT_US|UNSPECIFIED MONONEURITIS OF LOWER LIMB|UNSPECIFIED MONONEURITIS LOWER LIMB (DISORDER)
C0154747|T047|193154003|SNOMEDCT_US|MONONEURITIS LEG NOS|UNSPECIFIED MONONEURITIS LOWER LIMB (DISORDER)
C0154747|T047|193154003|SNOMEDCT_US|MONONEURITIS;LEGS|UNSPECIFIED MONONEURITIS LOWER LIMB (DISORDER)
C0154747|T047|193154003|SNOMEDCT_US|UNSPECIFIED MONONEURITIS LOWER LIMB |UNSPECIFIED MONONEURITIS LOWER LIMB (DISORDER)
C0154747|T047|193154003|SNOMEDCT_US|MONONEURITIS LOWER LIMB |UNSPECIFIED MONONEURITIS LOWER LIMB (DISORDER)
C0154747|T047|193154003|SNOMEDCT_US|UNSPECIFIED MONONEURITIS LOWER LIMB|UNSPECIFIED MONONEURITIS LOWER LIMB (DISORDER)
C0154747|T047|193154003|SNOMEDCT_US|MONONEURITIS OF LOWER LIMB |UNSPECIFIED MONONEURITIS LOWER LIMB (DISORDER)
C0154747|T047|193154003|SNOMEDCT_US|MONONEURITIS OF LOWER LIMB, UNSPECIFIED|UNSPECIFIED MONONEURITIS LOWER LIMB (DISORDER)
C0154747|T047|193154003|SNOMEDCT_US|LOWER LIMB; MONONEURITIS|UNSPECIFIED MONONEURITIS LOWER LIMB (DISORDER)
C0154747|T047|193154003|SNOMEDCT_US|MONONEURITIS; LOWER LIMB|UNSPECIFIED MONONEURITIS LOWER LIMB (DISORDER)
C0154747|T047|193154003|SNOMEDCT_US|MONONEURITIS OF LOWER LIMB, NOS|UNSPECIFIED MONONEURITIS LOWER LIMB (DISORDER)
C0154747|T047|193154003|SNOMEDCT_US|MONONEURITIS OF THE LEGS|UNSPECIFIED MONONEURITIS LOWER LIMB (DISORDER)
C0270890|T047|193123002|SNOMEDCT_US|NERVE ROOT AND PLEXUS DISORDERS|NERVE ROOT OR PLEXUS DISORDER NOS (DISORDER)
C0270890|T047|193123002|SNOMEDCT_US|NERVE ROOT AND PLEXUS DISORDER, UNSPECIFIED|NERVE ROOT OR PLEXUS DISORDER NOS (DISORDER)
C0270890|T047|193123002|SNOMEDCT_US|NERVE ROOT AND PLEXUS DISORDER |NERVE ROOT OR PLEXUS DISORDER NOS (DISORDER)
C0270890|T047|193123002|SNOMEDCT_US|NERVE ROOT AND PLEXUS DISORDER|NERVE ROOT OR PLEXUS DISORDER NOS (DISORDER)
C0270890|T047|193123002|SNOMEDCT_US|NERV ROOT/PLEXUS DIS NOS|NERVE ROOT OR PLEXUS DISORDER NOS (DISORDER)
C0270890|T047|193123002|SNOMEDCT_US|NERVE ROOT OR PLEXUS DISORDER NOS|NERVE ROOT OR PLEXUS DISORDER NOS (DISORDER)
C0270890|T047|193123002|SNOMEDCT_US|NERVE ROOT OR PLEXUS DISORDER NOS |NERVE ROOT OR PLEXUS DISORDER NOS (DISORDER)
C0270890|T047|193123002|SNOMEDCT_US|UNSPECIFIED NERVE ROOT AND PLEXUS DISORDER|NERVE ROOT OR PLEXUS DISORDER NOS (DISORDER)
C0270890|T047|193123002|SNOMEDCT_US|DISEASE (OR DISORDER); PLEXUS|NERVE ROOT OR PLEXUS DISORDER NOS (DISORDER)
C0435513|T047|208084009|SNOMEDCT_US|CLOSED FRACTURE OF COCCYX WITH COMPLETE CAUDA EQUINA LESION|CLOSED FRACTURE OF COCCYX WITH COMPLETE CAUDA EQUINA LESION (DISORDER)
C0435513|T047|208084009|SNOMEDCT_US|CLOSED FRACTURE OF COCCYX WITH COMPLETE CAUDA EQUINA LESION |CLOSED FRACTURE OF COCCYX WITH COMPLETE CAUDA EQUINA LESION (DISORDER)
C0435518|T047|208090008|SNOMEDCT_US|OPEN FRACTURE OF COCCYX WITH COMPLETE CAUDA EQUINA LESION|OPEN FRACTURE OF COCCYX WITH COMPLETE CAUDA EQUINA LESION (DISORDER)
C0435518|T047|208090008|SNOMEDCT_US|OPEN FRACTURE OF COCCYX WITH COMPLETE CAUDA EQUINA LESION |OPEN FRACTURE OF COCCYX WITH COMPLETE CAUDA EQUINA LESION (DISORDER)
C1960872|T047|426293000|SNOMEDCT_US|SURAL NEUROPATHY|SURAL NEUROPATHY (DISORDER)
C1960872|T047|426293000|SNOMEDCT_US|SURAL NEUROPATHY |SURAL NEUROPATHY (DISORDER)
C0435504|T047|208078006|SNOMEDCT_US|OPEN FRACTURE OF SACRUM WITH COMPLETE CAUDA EQUINA LESION|OPEN FRACTURE OF SACRUM WITH COMPLETE CAUDA EQUINA LESION (DISORDER)
C0435504|T047|208078006|SNOMEDCT_US|OPEN FRACTURE OF SACRUM WITH COMPLETE CAUDA EQUINA LESION |OPEN FRACTURE OF SACRUM WITH COMPLETE CAUDA EQUINA LESION (DISORDER)
C1268588|T047|129616004|SNOMEDCT_US|PORPHYRIC POLYNEUROPATHY|PORPHYRIC POLYNEUROPATHY (DISORDER)
C1268588|T047|129616004|SNOMEDCT_US|PORPHYRIC POLYNEUROPATHY |PORPHYRIC POLYNEUROPATHY (DISORDER)
C1268588|T047|129616004|SNOMEDCT_US|POLYNEUROPATHY IN PORPHYRIA |PORPHYRIC POLYNEUROPATHY (DISORDER)
C1268588|T047|129616004|SNOMEDCT_US|POLYNEUROPATHY IN PORPHYRIA|PORPHYRIC POLYNEUROPATHY (DISORDER)
C1268588|T047|129616004|SNOMEDCT_US|PORPHYRIC POLYNEUROPATHY |PORPHYRIC POLYNEUROPATHY (DISORDER)
C0032587|T047|128078004|SNOMEDCT_US|POLYRADICULONEUROPATHIES|POLYRADICULONEUROPATHY (DISORDER)
C0032587|T047|128078004|SNOMEDCT_US|POLYRADICULONEUROPATHY|POLYRADICULONEUROPATHY (DISORDER)
C0032587|T047|128078004|SNOMEDCT_US|POLYRADICULONEUROPATHY [DISEASE/FINDING]|POLYRADICULONEUROPATHY (DISORDER)
C0032587|T047|128078004|SNOMEDCT_US|POLYRADICULONEUROPATHY |POLYRADICULONEUROPATHY (DISORDER)
C0394023|T047|213197002|SNOMEDCT_US|DISRUPTION OF NERVE REPAIR|DISRUPTION OF NERVE REPAIR (DISORDER)
C0394023|T047|213197002|SNOMEDCT_US|DISRUPTION OF NERVE REPAIR |DISRUPTION OF NERVE REPAIR (DISORDER)
C0394025|T047|230805009|SNOMEDCT_US|NEUROMA OF NERVE REPAIR|NEUROMA OF NERVE REPAIR (DISORDER)
C0394025|T047|230805009|SNOMEDCT_US|NEUROMA OF NERVE REPAIR |NEUROMA OF NERVE REPAIR (DISORDER)
C0751929|T047|428461003|SNOMEDCT_US|NEUROPATHIES, SUPERFICIAL PERONEAL|SUPERFICIAL PERONEAL NERVE NEUROPATHY (DISORDER)
C0751929|T047|428461003|SNOMEDCT_US|PERONEAL NEUROPATHIES, SUPERFICIAL|SUPERFICIAL PERONEAL NERVE NEUROPATHY (DISORDER)
C0751929|T047|428461003|SNOMEDCT_US|PERONEAL NEUROPATHY, SUPERFICIAL|SUPERFICIAL PERONEAL NERVE NEUROPATHY (DISORDER)
C0751929|T047|428461003|SNOMEDCT_US|SUPERFICIAL PERONEAL NEUROPATHIES|SUPERFICIAL PERONEAL NERVE NEUROPATHY (DISORDER)
C0751929|T047|428461003|SNOMEDCT_US|SUPERFICIAL PERONEAL NEUROPATHY|SUPERFICIAL PERONEAL NERVE NEUROPATHY (DISORDER)
C0751929|T047|428461003|SNOMEDCT_US|SUPERFICIAL PERONEAL NERVE NEUROPATHY |SUPERFICIAL PERONEAL NERVE NEUROPATHY (DISORDER)
C0751929|T047|428461003|SNOMEDCT_US|SUPERFICIAL PERONEAL NERVE LESION|SUPERFICIAL PERONEAL NERVE NEUROPATHY (DISORDER)
C0751929|T047|428461003|SNOMEDCT_US|SUPERFICIAL PERONEAL NERVE NEUROPATHY|SUPERFICIAL PERONEAL NERVE NEUROPATHY (DISORDER)
C0751929|T047|428461003|SNOMEDCT_US|SUPERFICIAL PERONEAL NERVE DISORDER|SUPERFICIAL PERONEAL NERVE NEUROPATHY (DISORDER)
C0751929|T047|428461003|SNOMEDCT_US|SUPERFICIAL PERONEAL NERVE DISORDER |SUPERFICIAL PERONEAL NERVE NEUROPATHY (DISORDER)
C0751929|T047|428461003|SNOMEDCT_US|NEUROPATHY, SUPERFICIAL PERONEAL|SUPERFICIAL PERONEAL NERVE NEUROPATHY (DISORDER)
C2102996|T047||SNOMEDCT_US|DISORDERS OF PERIPHERAL NERVE, NEUROMUSCULAR JUNCTION AND MUSCLE 
C2102996|T047||SNOMEDCT_US|DISORDERS OF PERIPHERAL NERVE, NEUROMUSCULAR JUNCTION AND MUSCLE
C0442874|T047|386033004|SNOMEDCT_US|NEUROPATHY|NEUROPATHY (DISORDER)
C0442874|T047|386033004|SNOMEDCT_US|NERVE DISORDERS|NEUROPATHY (DISORDER)
C0442874|T047|386033004|SNOMEDCT_US|NERVE DISORDERS |NEUROPATHY (DISORDER)
C0442874|T047|386033004|SNOMEDCT_US|NEUROPATHY - (NOS)|NEUROPATHY (DISORDER)
C0442874|T047|386033004|SNOMEDCT_US|NEUROPATHY NOS|NEUROPATHY (DISORDER)
C0442874|T047|386033004|SNOMEDCT_US|NEUROPATHY |NEUROPATHY (DISORDER)
C0442874|T047|386033004|SNOMEDCT_US|NEUROPATHY (NERVE DAMAGE)|NEUROPATHY (DISORDER)
C0442874|T047|386033004|SNOMEDCT_US|NEUROPATHY |NEUROPATHY (DISORDER)
C0442874|T047|386033004|SNOMEDCT_US|NERVE; DISORDER|NEUROPATHY (DISORDER)
C0442874|T047|386033004|SNOMEDCT_US|NEUROPATHY, NOS|NEUROPATHY (DISORDER)
